* Library name: 6TSRAM_45n
* Cell name: bitcell_2X
* View name: schematic

.subckt bitcell_2X Q QB RBL RWL RWLB VDD VSS WBL WBLB WWL
 XM6 net1 QB VDD VDD pch_mac w=205.00n l=40n 
 XM5 net1 RWLB RBL VDD pch_mac w=205.00n l=40n
 XM4 Q QB VDD VDD pch_mac w=205.00n  l=40n
 XM3 QB Q VDD VDD pch_mac w=205.00n l=40n 
 XM9 WBL WWL Q VSS nch_mac w=310.0n  l=40n 
 XM8 WBLB WWL QB VSS nch_mac w=310.0n  l=40n 
 XM7 net1 QB VSS VSS nch_mac w=155.00n l=40n
 XM2 net1 RWL RBL VSS nch_mac w=155.00n  l=40n
 XM1 Q QB VSS VSS nch_mac w=155.00n l=40n
 XM0 QB Q VSS VSS nch_mac w=155.00n l=40n
.ends bitcell_2X
.SUBCKT array WWL3 WWL2 WWL1 WWL0 RWL3 RWL2 RWL1 RWL0 RWLB3
+ RWLB2 RWLB1 RWLB0 WBL15 WBL14 WBL13 WBL12 WBL11 WBL10
+ WBL9 WBL8 WBL7 WBL6 WBL5 WBL4 WBL3 WBL2 WBL1 WBL0
+ WBLB15 WBLB14 WBLB13 WBLB12 WBLB11 WBLB10 WBLB9 WBLB8 WBLB7
+ WBLB6 WBLB5 WBLB4 WBLB3 WBLB2 WBLB1 WBLB0 RBL15 RBL14
+ RBL13 RBL12 RBL11 RBL10 RBL9 RBL8 RBL7 RBL6 RBL5 RBL4
+ RBL3 RBL2 RBL1 RBL0 VDD VSS
    XI30 net0197 net0198 RBL5 RWL1 RWLB1 VDD VSS WBL5 WBLB5 WWL1 \
        bitcell_2X
    XI33 net0191 net0192 RBL4 RWL0 RWLB0 VDD VSS WBL4 WBLB4 WWL0 \
        bitcell_2X
    XI17 net0223 net0224 RBL2 RWL1 RWLB1 VDD VSS WBL2 WBLB2 WWL1 \
        bitcell_2X
    XI42 net0173 net0174 RBL9 RWL3 RWLB3 VDD VSS WBL9 WBLB9 WWL3 \
        bitcell_2X
    XI26 net0205 net0206 RBL4 RWL2 RWLB2 VDD VSS WBL4 WBLB4 WWL2 \
        bitcell_2X
    XI67 net0123 net0124 RBL11 RWL0 RWLB0 VDD VSS WBL11 WBLB11 WWL0 \
        bitcell_2X
    XI11 net0235 net0236 RBL1 RWL2 RWLB2 VDD VSS WBL1 WBLB1 WWL2 \
        bitcell_2X
    XI50 net0157 net0158 RBL14 RWL1 RWLB1 VDD VSS WBL14 WBLB14 WWL1 \
        bitcell_2X
    XI27 net0203 net0204 RBL6 RWL2 RWLB2 VDD VSS WBL6 WBLB6 WWL2 \
        bitcell_2X
    XI34 net0189 net0190 RBL5 RWL0 RWLB0 VDD VSS WBL5 WBLB5 WWL0 \
        bitcell_2X
    XI18 net0221 net0222 RBL3 RWL1 RWLB1 VDD VSS WBL3 WBLB3 WWL1 \
        bitcell_2X
    XI61 net0135 net0136 RBL8 RWL1 RWLB1 VDD VSS WBL8 WBLB8 WWL1 \
        bitcell_2X
    XI35 net0187 net0188 RBL7 RWL0 RWLB0 VDD VSS WBL7 WBLB7 WWL0 \
        bitcell_2X
    XI43 net0171 net0172 RBL11 RWL3 RWLB3 VDD VSS WBL11 WBLB11 WWL3 \
        bitcell_2X
    XI19 net0219 net0220 RBL2 RWL0 RWLB0 VDD VSS WBL2 WBLB2 WWL0 \
        bitcell_2X
    XI28 net0201 net0202 RBL7 RWL2 RWLB2 VDD VSS WBL7 WBLB7 WWL2 \
        bitcell_2X
    XI44 net0169 net0170 RBL10 RWL3 RWLB3 VDD VSS WBL10 WBLB10 WWL3 \
        bitcell_2X
    XI68 net0121 net0122 RBL10 RWL0 RWLB0 VDD VSS WBL10 WBLB10 WWL0 \
        bitcell_2X
    XI51 net0155 net0156 RBL15 RWL1 RWLB1 VDD VSS WBL15 WBLB15 WWL1 \
        bitcell_2X
    XI12 net0233 net0234 RBL1 RWL0 RWLB0 VDD VSS WBL1 WBLB1 WWL0 \
        bitcell_2X
    XI62 net0133 net0134 RBL9 RWL1 RWLB1 VDD VSS WBL9 WBLB9 WWL1 \
        bitcell_2X
    XI36 net0185 net0186 RBL6 RWL0 RWLB0 VDD VSS WBL6 WBLB6 WWL0 \
        bitcell_2X
    XI29 net0199 net0200 RBL4 RWL1 RWLB1 VDD VSS WBL4 WBLB4 WWL1 \
        bitcell_2X
    XI20 net0217 net0218 RBL3 RWL0 RWLB0 VDD VSS WBL3 WBLB3 WWL0 \
        bitcell_2X
    XI45 net0167 net0168 RBL13 RWL2 RWLB2 VDD VSS WBL13 WBLB13 WWL2 \
        bitcell_2X
    XI63 net0131 net0132 RBL11 RWL1 RWLB1 VDD VSS WBL11 WBLB11 WWL1 \
        bitcell_2X
    XI52 net0153 net0154 RBL13 RWL1 RWLB1 VDD VSS WBL13 WBLB13 WWL1 \
        bitcell_2X
    XI37 net0183 net0184 RBL8 RWL3 RWLB3 VDD VSS WBL8 WBLB8 WWL3 \
        bitcell_2X
    XI13 net0231 net0232 RBL2 RWL3 RWLB3 VDD VSS WBL2 WBLB2 WWL3 \
        bitcell_2X
    XI53 net0151 net0152 RBL12 RWL1 RWLB1 VDD VSS WBL12 WBLB12 WWL1 \
        bitcell_2X
    XI14 net0229 net0230 RBL3 RWL3 RWLB3 VDD VSS WBL3 WBLB3 WWL3 \
        bitcell_2X
    XI38 net0181 net0182 RBL15 RWL3 RWLB3 VDD VSS WBL15 WBLB15 WWL3 \
        bitcell_2X
    XI66 net0125 net0126 RBL9 RWL0 RWLB0 VDD VSS WBL9 WBLB9 WWL0 \
        bitcell_2X
    XI65 net0127 net0128 RBL8 RWL0 RWLB0 VDD VSS WBL8 WBLB8 WWL0 \
        bitcell_2X
    XI48 net0161 net0162 RBL13 RWL0 RWLB0 VDD VSS WBL13 WBLB13 WWL0 \
        bitcell_2X
    XI46 net0165 net0166 RBL14 RWL0 RWLB0 VDD VSS WBL14 WBLB14 WWL0 \
        bitcell_2X
    XI9 net0239 net0240 RBL1 RWL3 RWLB3 VDD VSS WBL1 WBLB1 WWL3 \
        bitcell_2X
    XI58 net0141 net0142 RBL8 RWL2 RWLB2 VDD VSS WBL8 WBLB8 WWL2 \
        bitcell_2X
    XI39 net0179 net0180 RBL14 RWL3 RWLB3 VDD VSS WBL14 WBLB14 WWL3 \
        bitcell_2X
    XI6 net20 net21 RBL0 RWL1 RWLB1 VDD VSS WBL0 WBLB0 WWL1 bitcell_2X
    XI10 net0237 net0238 RBL1 RWL1 RWLB1 VDD VSS WBL1 WBLB1 WWL1 \
        bitcell_2X
    XI59 net0139 net0140 RBL10 RWL2 RWLB2 VDD VSS WBL10 WBLB10 WWL2 \
        bitcell_2X
    XI40 net0177 net0178 RBL12 RWL3 RWLB3 VDD VSS WBL12 WBLB12 WWL3 \
        bitcell_2X
    XI22 net0213 net0214 RBL5 RWL3 RWLB3 VDD VSS WBL5 WBLB5 WWL3 \
        bitcell_2X
    XI21 net0215 net0216 RBL4 RWL3 RWLB3 VDD VSS WBL4 WBLB4 WWL3 \
        bitcell_2X
    XI56 net0145 net0146 RBL12 RWL2 RWLB2 VDD VSS WBL12 WBLB12 WWL2 \
        bitcell_2X
    XI32 net0193 net0194 RBL6 RWL1 RWLB1 VDD VSS WBL6 WBLB6 WWL1 \
        bitcell_2X
    XI47 net0163 net0164 RBL15 RWL0 RWLB0 VDD VSS WBL15 WBLB15 WWL0 \
        bitcell_2X
    XI64 net0129 net0130 RBL10 RWL1 RWLB1 VDD VSS WBL10 WBLB10 WWL1 \
        bitcell_2X
    XI57 net0143 net0144 RBL9 RWL2 RWLB2 VDD VSS WBL9 WBLB9 WWL2 \
        bitcell_2X
    XI55 net0147 net0148 RBL14 RWL2 RWLB2 VDD VSS WBL14 WBLB14 WWL2 \
        bitcell_2X
    XI54 net0149 net0150 RBL15 RWL2 RWLB2 VDD VSS WBL15 WBLB15 WWL2 \
        bitcell_2X
    XI49 net0159 net0160 RBL12 RWL0 RWLB0 VDD VSS WBL12 WBLB12 WWL0 \
        bitcell_2X
    XI16 net0225 net0226 RBL2 RWL2 RWLB2 VDD VSS WBL2 WBLB2 WWL2 \
        bitcell_2X
    XI31 net0195 net0196 RBL7 RWL1 RWLB1 VDD VSS WBL7 WBLB7 WWL1 \
        bitcell_2X
    XI15 net0227 net0228 RBL3 RWL2 RWLB2 VDD VSS WBL3 WBLB3 WWL2 \
        bitcell_2X
    XI60 net0137 net0138 RBL11 RWL2 RWLB2 VDD VSS WBL11 WBLB11 WWL2 \
        bitcell_2X
    XI41 net0175 net0176 RBL13 RWL3 RWLB3 VDD VSS WBL13 WBLB13 WWL3 \
        bitcell_2X
    XI24 net0209 net0210 RBL6 RWL3 RWLB3 VDD VSS WBL6 WBLB6 WWL3 \
        bitcell_2X
    XI7 net18 net19 RBL0 RWL2 RWLB2 VDD VSS WBL0 WBLB0 WWL2 bitcell_2X
    XI23 net0211 net0212 RBL7 RWL3 RWLB3 VDD VSS WBL7 WBLB7 WWL3 \
        bitcell_2X
    XI4 net22 net23 RBL0 RWL0 RWLB0 VDD VSS WBL0 WBLB0 WWL0 bitcell_2X
    XI25 net0207 net0208 RBL5 RWL2 RWLB2 VDD VSS WBL5 WBLB5 WWL2 \
        bitcell_2X
    XI8 net16 net17 RBL0 RWL3 RWLB3 VDD VSS WBL0 WBLB0 WWL3 bitcell_2X
.ends array

