************************************************************************
* auCdl Netlist:
* 
* Library Name:  10T
* Top Cell Name: 16x16_10T_new
* View Name:     schematic
* Netlisted on:  Aug  9 09:09:14 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: 10T
* Cell Name:    10TSRAM_M8
* View Name:    schematic
************************************************************************

.SUBCKT 10TSRAM_M8 GND RBL RWL RWLB VDD WBL WBLB WWLB
*.PININFO GND:I RWL:I RWLB:I VDD:I WBL:I WBLB:I WWLB:I RBL:O
MM8 net08 RWL RBL GND nch l=60n w=120.0n m=1
MM7 net08 QB GND GND nch l=60n w=160.0n m=1
MM10 WBL WWLB Q GND nch l=60n w=180.0n m=1
MM11 WBLB WWLB QB GND nch l=60n w=180.0n m=1
MM1 Q QB GND GND nch l=60n w=120.0n m=1
MM0 QB Q GND GND nch l=60n w=120.0n m=1
MM9 net08 RWLB RBL VDD pch l=60n w=120.0n m=1
MM6 net08 QB VDD VDD pch l=60n w=480.0n m=1
MM5 Q QB VDD VDD pch l=60n w=240.0n m=1
MM4 QB Q VDD VDD pch l=60n w=240.0n m=1
.ENDS

************************************************************************
* Library Name: 10T
* Cell Name:    16x16_10T_new
* View Name:    schematic
************************************************************************

.SUBCKT array GND RBL[0] RBL[1] RBL[2] RBL[3] RBL[4] RBL[5] RBL[6] 
+ RBL[7] RBL[8] RBL[9] RBL[10] RBL[11] RBL[12] RBL[13] RBL[14] RBL[15] RWL[0] 
+ RWL[1] RWL[2] RWL[3] RWL[4] RWL[5] RWL[6] RWL[7] RWL[8] RWL[9] RWL[10] 
+ RWL[11] RWL[12] RWL[13] RWL[14] RWL[15] RWLB[0] RWLB[1] RWLB[2] RWLB[3] 
+ RWLB[4] RWLB[5] RWLB[6] RWLB[7] RWLB[8] RWLB[9] RWLB[10] RWLB[11] RWLB[12] 
+ RWLB[13] RWLB[14] RWLB[15] VDD WBL[0] WBL[1] WBL[2] WBL[3] WBL[4] WBL[5] 
+ WBL[6] WBL[7] WBL[8] WBL[9] WBL[10] WBL[11] WBL[12] WBL[13] WBL[14] WBL[15] 
+ WBLB[0] WBLB[1] WBLB[2] WBLB[3] WBLB[4] WBLB[5] WBLB[6] WBLB[7] WBLB[8] 
+ WBLB[9] WBLB[10] WBLB[11] WBLB[12] WBLB[13] WBLB[14] WBLB[15] WWLB[0] 
+ WWLB[1] WWLB[2] WWLB[3] WWLB[4] WWLB[5] WWLB[6] WWLB[7] WWLB[8] WWLB[9] 
+ WWLB[10] WWLB[11] WWLB[12] WWLB[13] WWLB[14] WWLB[15]
*.PININFO RWL[0]:I RWL[1]:I RWL[2]:I RWL[3]:I RWL[4]:I RWL[5]:I RWL[6]:I 
*.PININFO RWL[7]:I RWL[8]:I RWL[9]:I RWL[10]:I RWL[11]:I RWL[12]:I RWL[13]:I 
*.PININFO RWL[14]:I RWL[15]:I RWLB[0]:I RWLB[1]:I RWLB[2]:I RWLB[3]:I 
*.PININFO RWLB[4]:I RWLB[5]:I RWLB[6]:I RWLB[7]:I RWLB[8]:I RWLB[9]:I 
*.PININFO RWLB[10]:I RWLB[11]:I RWLB[12]:I RWLB[13]:I RWLB[14]:I RWLB[15]:I 
*.PININFO WBL[0]:I WBL[1]:I WBL[2]:I WBL[3]:I WBL[4]:I WBL[5]:I WBL[6]:I 
*.PININFO WBL[7]:I WBL[8]:I WBL[9]:I WBL[10]:I WBL[11]:I WBL[12]:I WBL[13]:I 
*.PININFO WBL[14]:I WBL[15]:I WBLB[0]:I WBLB[1]:I WBLB[2]:I WBLB[3]:I 
*.PININFO WBLB[4]:I WBLB[5]:I WBLB[6]:I WBLB[7]:I WBLB[8]:I WBLB[9]:I 
*.PININFO WBLB[10]:I WBLB[11]:I WBLB[12]:I WBLB[13]:I WBLB[14]:I WBLB[15]:I 
*.PININFO WWLB[0]:I WWLB[1]:I WWLB[2]:I WWLB[3]:I WWLB[4]:I WWLB[5]:I 
*.PININFO WWLB[6]:I WWLB[7]:I WWLB[8]:I WWLB[9]:I WWLB[10]:I WWLB[11]:I 
*.PININFO WWLB[12]:I WWLB[13]:I WWLB[14]:I WWLB[15]:I RBL[0]:O RBL[1]:O 
*.PININFO RBL[2]:O RBL[3]:O RBL[4]:O RBL[5]:O RBL[6]:O RBL[7]:O RBL[8]:O 
*.PININFO RBL[9]:O RBL[10]:O RBL[11]:O RBL[12]:O RBL[13]:O RBL[14]:O RBL[15]:O 
*.PININFO GND:B VDD:B
XI1006 GND RBL[14] RWL[14] RWLB[14] VDD WBL[14] WBLB[14] WWLB[14] / 10TSRAM_M8
XI1020 GND RBL[0] RWL[14] RWLB[14] VDD WBL[0] WBLB[0] WWLB[14] / 10TSRAM_M8
XI1019 GND RBL[1] RWL[14] RWLB[14] VDD WBL[1] WBLB[1] WWLB[14] / 10TSRAM_M8
XI1018 GND RBL[2] RWL[14] RWLB[14] VDD WBL[2] WBLB[2] WWLB[14] / 10TSRAM_M8
XI1017 GND RBL[3] RWL[14] RWLB[14] VDD WBL[3] WBLB[3] WWLB[14] / 10TSRAM_M8
XI1016 GND RBL[4] RWL[14] RWLB[14] VDD WBL[4] WBLB[4] WWLB[14] / 10TSRAM_M8
XI1015 GND RBL[5] RWL[14] RWLB[14] VDD WBL[5] WBLB[5] WWLB[14] / 10TSRAM_M8
XI1014 GND RBL[6] RWL[14] RWLB[14] VDD WBL[6] WBLB[6] WWLB[14] / 10TSRAM_M8
XI1013 GND RBL[7] RWL[14] RWLB[14] VDD WBL[7] WBLB[7] WWLB[14] / 10TSRAM_M8
XI1012 GND RBL[8] RWL[14] RWLB[14] VDD WBL[8] WBLB[8] WWLB[14] / 10TSRAM_M8
XI1011 GND RBL[9] RWL[14] RWLB[14] VDD WBL[9] WBLB[9] WWLB[14] / 10TSRAM_M8
XI1010 GND RBL[10] RWL[14] RWLB[14] VDD WBL[10] WBLB[10] WWLB[14] / 10TSRAM_M8
XI1009 GND RBL[11] RWL[14] RWLB[14] VDD WBL[11] WBLB[11] WWLB[14] / 10TSRAM_M8
XI1008 GND RBL[12] RWL[14] RWLB[14] VDD WBL[12] WBLB[12] WWLB[14] / 10TSRAM_M8
XI1007 GND RBL[13] RWL[14] RWLB[14] VDD WBL[13] WBLB[13] WWLB[14] / 10TSRAM_M8
XI1021 GND RBL[15] RWL[14] RWLB[14] VDD WBL[15] WBLB[15] WWLB[14] / 10TSRAM_M8
XI1037 GND RBL[15] RWL[15] RWLB[15] VDD WBL[15] WBLB[15] WWLB[15] / 10TSRAM_M8
XI1036 GND RBL[0] RWL[15] RWLB[15] VDD WBL[0] WBLB[0] WWLB[15] / 10TSRAM_M8
XI984 GND RBL[4] RWL[12] RWLB[12] VDD WBL[4] WBLB[4] WWLB[12] / 10TSRAM_M8
XI1035 GND RBL[1] RWL[15] RWLB[15] VDD WBL[1] WBLB[1] WWLB[15] / 10TSRAM_M8
XI992 GND RBL[12] RWL[13] RWLB[13] VDD WBL[12] WBLB[12] WWLB[13] / 10TSRAM_M8
XI951 GND RBL[5] RWL[10] RWLB[10] VDD WBL[5] WBLB[5] WWLB[10] / 10TSRAM_M8
XI950 GND RBL[6] RWL[10] RWLB[10] VDD WBL[6] WBLB[6] WWLB[10] / 10TSRAM_M8
XI949 GND RBL[7] RWL[10] RWLB[10] VDD WBL[7] WBLB[7] WWLB[10] / 10TSRAM_M8
XI948 GND RBL[8] RWL[10] RWLB[10] VDD WBL[8] WBLB[8] WWLB[10] / 10TSRAM_M8
XI975 GND RBL[13] RWL[12] RWLB[12] VDD WBL[13] WBLB[13] WWLB[12] / 10TSRAM_M8
XI974 GND RBL[14] RWL[12] RWLB[12] VDD WBL[14] WBLB[14] WWLB[12] / 10TSRAM_M8
XI973 GND RBL[15] RWL[11] RWLB[11] VDD WBL[15] WBLB[15] WWLB[11] / 10TSRAM_M8
XI972 GND RBL[0] RWL[11] RWLB[11] VDD WBL[0] WBLB[0] WWLB[11] / 10TSRAM_M8
XI971 GND RBL[1] RWL[11] RWLB[11] VDD WBL[1] WBLB[1] WWLB[11] / 10TSRAM_M8
XI970 GND RBL[2] RWL[11] RWLB[11] VDD WBL[2] WBLB[2] WWLB[11] / 10TSRAM_M8
XI990 GND RBL[14] RWL[13] RWLB[13] VDD WBL[14] WBLB[14] WWLB[13] / 10TSRAM_M8
XI989 GND RBL[15] RWL[12] RWLB[12] VDD WBL[15] WBLB[15] WWLB[12] / 10TSRAM_M8
XI988 GND RBL[0] RWL[12] RWLB[12] VDD WBL[0] WBLB[0] WWLB[12] / 10TSRAM_M8
XI991 GND RBL[13] RWL[13] RWLB[13] VDD WBL[13] WBLB[13] WWLB[13] / 10TSRAM_M8
XI981 GND RBL[7] RWL[12] RWLB[12] VDD WBL[7] WBLB[7] WWLB[12] / 10TSRAM_M8
XI980 GND RBL[8] RWL[12] RWLB[12] VDD WBL[8] WBLB[8] WWLB[12] / 10TSRAM_M8
XI1034 GND RBL[2] RWL[15] RWLB[15] VDD WBL[2] WBLB[2] WWLB[15] / 10TSRAM_M8
XI993 GND RBL[11] RWL[13] RWLB[13] VDD WBL[11] WBLB[11] WWLB[13] / 10TSRAM_M8
XI947 GND RBL[9] RWL[10] RWLB[10] VDD WBL[9] WBLB[9] WWLB[10] / 10TSRAM_M8
XI946 GND RBL[10] RWL[10] RWLB[10] VDD WBL[10] WBLB[10] WWLB[10] / 10TSRAM_M8
XI945 GND RBL[11] RWL[10] RWLB[10] VDD WBL[11] WBLB[11] WWLB[10] / 10TSRAM_M8
XI944 GND RBL[12] RWL[10] RWLB[10] VDD WBL[12] WBLB[12] WWLB[10] / 10TSRAM_M8
XI969 GND RBL[3] RWL[11] RWLB[11] VDD WBL[3] WBLB[3] WWLB[11] / 10TSRAM_M8
XI968 GND RBL[4] RWL[11] RWLB[11] VDD WBL[4] WBLB[4] WWLB[11] / 10TSRAM_M8
XI967 GND RBL[5] RWL[11] RWLB[11] VDD WBL[5] WBLB[5] WWLB[11] / 10TSRAM_M8
XI966 GND RBL[6] RWL[11] RWLB[11] VDD WBL[6] WBLB[6] WWLB[11] / 10TSRAM_M8
XI965 GND RBL[7] RWL[11] RWLB[11] VDD WBL[7] WBLB[7] WWLB[11] / 10TSRAM_M8
XI964 GND RBL[8] RWL[11] RWLB[11] VDD WBL[8] WBLB[8] WWLB[11] / 10TSRAM_M8
XI987 GND RBL[1] RWL[12] RWLB[12] VDD WBL[1] WBLB[1] WWLB[12] / 10TSRAM_M8
XI986 GND RBL[2] RWL[12] RWLB[12] VDD WBL[2] WBLB[2] WWLB[12] / 10TSRAM_M8
XI985 GND RBL[3] RWL[12] RWLB[12] VDD WBL[3] WBLB[3] WWLB[12] / 10TSRAM_M8
XI978 GND RBL[10] RWL[12] RWLB[12] VDD WBL[10] WBLB[10] WWLB[12] / 10TSRAM_M8
XI977 GND RBL[11] RWL[12] RWLB[12] VDD WBL[11] WBLB[11] WWLB[12] / 10TSRAM_M8
XI976 GND RBL[12] RWL[12] RWLB[12] VDD WBL[12] WBLB[12] WWLB[12] / 10TSRAM_M8
XI1033 GND RBL[3] RWL[15] RWLB[15] VDD WBL[3] WBLB[3] WWLB[15] / 10TSRAM_M8
XI994 GND RBL[10] RWL[13] RWLB[13] VDD WBL[10] WBLB[10] WWLB[13] / 10TSRAM_M8
XI943 GND RBL[13] RWL[10] RWLB[10] VDD WBL[13] WBLB[13] WWLB[10] / 10TSRAM_M8
XI942 GND RBL[14] RWL[10] RWLB[10] VDD WBL[14] WBLB[14] WWLB[10] / 10TSRAM_M8
XI941 GND RBL[15] RWL[9] RWLB[9] VDD WBL[15] WBLB[15] WWLB[9] / 10TSRAM_M8
XI940 GND RBL[0] RWL[9] RWLB[9] VDD WBL[0] WBLB[0] WWLB[9] / 10TSRAM_M8
XI963 GND RBL[9] RWL[11] RWLB[11] VDD WBL[9] WBLB[9] WWLB[11] / 10TSRAM_M8
XI962 GND RBL[10] RWL[11] RWLB[11] VDD WBL[10] WBLB[10] WWLB[11] / 10TSRAM_M8
XI961 GND RBL[11] RWL[11] RWLB[11] VDD WBL[11] WBLB[11] WWLB[11] / 10TSRAM_M8
XI960 GND RBL[12] RWL[11] RWLB[11] VDD WBL[12] WBLB[12] WWLB[11] / 10TSRAM_M8
XI959 GND RBL[13] RWL[11] RWLB[11] VDD WBL[13] WBLB[13] WWLB[11] / 10TSRAM_M8
XI958 GND RBL[14] RWL[11] RWLB[11] VDD WBL[14] WBLB[14] WWLB[11] / 10TSRAM_M8
XI983 GND RBL[5] RWL[12] RWLB[12] VDD WBL[5] WBLB[5] WWLB[12] / 10TSRAM_M8
XI982 GND RBL[6] RWL[12] RWLB[12] VDD WBL[6] WBLB[6] WWLB[12] / 10TSRAM_M8
XI934 GND RBL[6] RWL[9] RWLB[9] VDD WBL[6] WBLB[6] WWLB[9] / 10TSRAM_M8
XI933 GND RBL[7] RWL[9] RWLB[9] VDD WBL[7] WBLB[7] WWLB[9] / 10TSRAM_M8
XI932 GND RBL[8] RWL[9] RWLB[9] VDD WBL[8] WBLB[8] WWLB[9] / 10TSRAM_M8
XI935 GND RBL[5] RWL[9] RWLB[9] VDD WBL[5] WBLB[5] WWLB[9] / 10TSRAM_M8
XI1032 GND RBL[4] RWL[15] RWLB[15] VDD WBL[4] WBLB[4] WWLB[15] / 10TSRAM_M8
XI995 GND RBL[9] RWL[13] RWLB[13] VDD WBL[9] WBLB[9] WWLB[13] / 10TSRAM_M8
XI938 GND RBL[2] RWL[9] RWLB[9] VDD WBL[2] WBLB[2] WWLB[9] / 10TSRAM_M8
XI937 GND RBL[3] RWL[9] RWLB[9] VDD WBL[3] WBLB[3] WWLB[9] / 10TSRAM_M8
XI936 GND RBL[4] RWL[9] RWLB[9] VDD WBL[4] WBLB[4] WWLB[9] / 10TSRAM_M8
XI939 GND RBL[1] RWL[9] RWLB[9] VDD WBL[1] WBLB[1] WWLB[9] / 10TSRAM_M8
XI956 GND RBL[0] RWL[10] RWLB[10] VDD WBL[0] WBLB[0] WWLB[10] / 10TSRAM_M8
XI955 GND RBL[1] RWL[10] RWLB[10] VDD WBL[1] WBLB[1] WWLB[10] / 10TSRAM_M8
XI954 GND RBL[2] RWL[10] RWLB[10] VDD WBL[2] WBLB[2] WWLB[10] / 10TSRAM_M8
XI953 GND RBL[3] RWL[10] RWLB[10] VDD WBL[3] WBLB[3] WWLB[10] / 10TSRAM_M8
XI952 GND RBL[4] RWL[10] RWLB[10] VDD WBL[4] WBLB[4] WWLB[10] / 10TSRAM_M8
XI957 GND RBL[15] RWL[10] RWLB[10] VDD WBL[15] WBLB[15] WWLB[10] / 10TSRAM_M8
XI979 GND RBL[9] RWL[12] RWLB[12] VDD WBL[9] WBLB[9] WWLB[12] / 10TSRAM_M8
XI900 GND RBL[8] RWL[7] RWLB[7] VDD WBL[8] WBLB[8] WWLB[7] / 10TSRAM_M8
XI931 GND RBL[9] RWL[9] RWLB[9] VDD WBL[9] WBLB[9] WWLB[9] / 10TSRAM_M8
XI930 GND RBL[10] RWL[9] RWLB[9] VDD WBL[10] WBLB[10] WWLB[9] / 10TSRAM_M8
XI929 GND RBL[11] RWL[9] RWLB[9] VDD WBL[11] WBLB[11] WWLB[9] / 10TSRAM_M8
XI928 GND RBL[12] RWL[9] RWLB[9] VDD WBL[12] WBLB[12] WWLB[9] / 10TSRAM_M8
XI1031 GND RBL[5] RWL[15] RWLB[15] VDD WBL[5] WBLB[5] WWLB[15] / 10TSRAM_M8
XI996 GND RBL[8] RWL[13] RWLB[13] VDD WBL[8] WBLB[8] WWLB[13] / 10TSRAM_M8
XI875 GND RBL[1] RWL[5] RWLB[5] VDD WBL[1] WBLB[1] WWLB[5] / 10TSRAM_M8
XI874 GND RBL[2] RWL[5] RWLB[5] VDD WBL[2] WBLB[2] WWLB[5] / 10TSRAM_M8
XI873 GND RBL[3] RWL[5] RWLB[5] VDD WBL[3] WBLB[3] WWLB[5] / 10TSRAM_M8
XI872 GND RBL[4] RWL[5] RWLB[5] VDD WBL[4] WBLB[4] WWLB[5] / 10TSRAM_M8
XI911 GND RBL[13] RWL[8] RWLB[8] VDD WBL[13] WBLB[13] WWLB[8] / 10TSRAM_M8
XI910 GND RBL[14] RWL[8] RWLB[8] VDD WBL[14] WBLB[14] WWLB[8] / 10TSRAM_M8
XI909 GND RBL[15] RWL[7] RWLB[7] VDD WBL[15] WBLB[15] WWLB[7] / 10TSRAM_M8
XI908 GND RBL[0] RWL[7] RWLB[7] VDD WBL[0] WBLB[0] WWLB[7] / 10TSRAM_M8
XI907 GND RBL[1] RWL[7] RWLB[7] VDD WBL[1] WBLB[1] WWLB[7] / 10TSRAM_M8
XI906 GND RBL[2] RWL[7] RWLB[7] VDD WBL[2] WBLB[2] WWLB[7] / 10TSRAM_M8
XI895 GND RBL[13] RWL[7] RWLB[7] VDD WBL[13] WBLB[13] WWLB[7] / 10TSRAM_M8
XI894 GND RBL[14] RWL[7] RWLB[7] VDD WBL[14] WBLB[14] WWLB[7] / 10TSRAM_M8
XI927 GND RBL[13] RWL[9] RWLB[9] VDD WBL[13] WBLB[13] WWLB[9] / 10TSRAM_M8
XI926 GND RBL[14] RWL[9] RWLB[9] VDD WBL[14] WBLB[14] WWLB[9] / 10TSRAM_M8
XI925 GND RBL[15] RWL[8] RWLB[8] VDD WBL[15] WBLB[15] WWLB[8] / 10TSRAM_M8
XI924 GND RBL[0] RWL[8] RWLB[8] VDD WBL[0] WBLB[0] WWLB[8] / 10TSRAM_M8
XI1030 GND RBL[6] RWL[15] RWLB[15] VDD WBL[6] WBLB[6] WWLB[15] / 10TSRAM_M8
XI997 GND RBL[7] RWL[13] RWLB[13] VDD WBL[7] WBLB[7] WWLB[13] / 10TSRAM_M8
XI871 GND RBL[5] RWL[5] RWLB[5] VDD WBL[5] WBLB[5] WWLB[5] / 10TSRAM_M8
XI870 GND RBL[6] RWL[5] RWLB[5] VDD WBL[6] WBLB[6] WWLB[5] / 10TSRAM_M8
XI869 GND RBL[7] RWL[5] RWLB[5] VDD WBL[7] WBLB[7] WWLB[5] / 10TSRAM_M8
XI868 GND RBL[8] RWL[5] RWLB[5] VDD WBL[8] WBLB[8] WWLB[5] / 10TSRAM_M8
XI905 GND RBL[3] RWL[7] RWLB[7] VDD WBL[3] WBLB[3] WWLB[7] / 10TSRAM_M8
XI904 GND RBL[4] RWL[7] RWLB[7] VDD WBL[4] WBLB[4] WWLB[7] / 10TSRAM_M8
XI903 GND RBL[5] RWL[7] RWLB[7] VDD WBL[5] WBLB[5] WWLB[7] / 10TSRAM_M8
XI902 GND RBL[6] RWL[7] RWLB[7] VDD WBL[6] WBLB[6] WWLB[7] / 10TSRAM_M8
XI901 GND RBL[7] RWL[7] RWLB[7] VDD WBL[7] WBLB[7] WWLB[7] / 10TSRAM_M8
XI890 GND RBL[2] RWL[6] RWLB[6] VDD WBL[2] WBLB[2] WWLB[6] / 10TSRAM_M8
XI889 GND RBL[3] RWL[6] RWLB[6] VDD WBL[3] WBLB[3] WWLB[6] / 10TSRAM_M8
XI888 GND RBL[4] RWL[6] RWLB[6] VDD WBL[4] WBLB[4] WWLB[6] / 10TSRAM_M8
XI923 GND RBL[1] RWL[8] RWLB[8] VDD WBL[1] WBLB[1] WWLB[8] / 10TSRAM_M8
XI922 GND RBL[2] RWL[8] RWLB[8] VDD WBL[2] WBLB[2] WWLB[8] / 10TSRAM_M8
XI921 GND RBL[3] RWL[8] RWLB[8] VDD WBL[3] WBLB[3] WWLB[8] / 10TSRAM_M8
XI920 GND RBL[4] RWL[8] RWLB[8] VDD WBL[4] WBLB[4] WWLB[8] / 10TSRAM_M8
XI1029 GND RBL[7] RWL[15] RWLB[15] VDD WBL[7] WBLB[7] WWLB[15] / 10TSRAM_M8
XI998 GND RBL[6] RWL[13] RWLB[13] VDD WBL[6] WBLB[6] WWLB[13] / 10TSRAM_M8
XI867 GND RBL[9] RWL[5] RWLB[5] VDD WBL[9] WBLB[9] WWLB[5] / 10TSRAM_M8
XI866 GND RBL[10] RWL[5] RWLB[5] VDD WBL[10] WBLB[10] WWLB[5] / 10TSRAM_M8
XI865 GND RBL[11] RWL[5] RWLB[5] VDD WBL[11] WBLB[11] WWLB[5] / 10TSRAM_M8
XI864 GND RBL[12] RWL[5] RWLB[5] VDD WBL[12] WBLB[12] WWLB[5] / 10TSRAM_M8
XI899 GND RBL[9] RWL[7] RWLB[7] VDD WBL[9] WBLB[9] WWLB[7] / 10TSRAM_M8
XI898 GND RBL[10] RWL[7] RWLB[7] VDD WBL[10] WBLB[10] WWLB[7] / 10TSRAM_M8
XI897 GND RBL[11] RWL[7] RWLB[7] VDD WBL[11] WBLB[11] WWLB[7] / 10TSRAM_M8
XI896 GND RBL[12] RWL[7] RWLB[7] VDD WBL[12] WBLB[12] WWLB[7] / 10TSRAM_M8
XI885 GND RBL[7] RWL[6] RWLB[6] VDD WBL[7] WBLB[7] WWLB[6] / 10TSRAM_M8
XI884 GND RBL[8] RWL[6] RWLB[6] VDD WBL[8] WBLB[8] WWLB[6] / 10TSRAM_M8
XI883 GND RBL[9] RWL[6] RWLB[6] VDD WBL[9] WBLB[9] WWLB[6] / 10TSRAM_M8
XI882 GND RBL[10] RWL[6] RWLB[6] VDD WBL[10] WBLB[10] WWLB[6] / 10TSRAM_M8
XI919 GND RBL[5] RWL[8] RWLB[8] VDD WBL[5] WBLB[5] WWLB[8] / 10TSRAM_M8
XI918 GND RBL[6] RWL[8] RWLB[8] VDD WBL[6] WBLB[6] WWLB[8] / 10TSRAM_M8
XI917 GND RBL[7] RWL[8] RWLB[8] VDD WBL[7] WBLB[7] WWLB[8] / 10TSRAM_M8
XI916 GND RBL[8] RWL[8] RWLB[8] VDD WBL[8] WBLB[8] WWLB[8] / 10TSRAM_M8
XI1028 GND RBL[8] RWL[15] RWLB[15] VDD WBL[8] WBLB[8] WWLB[15] / 10TSRAM_M8
XI999 GND RBL[5] RWL[13] RWLB[13] VDD WBL[5] WBLB[5] WWLB[13] / 10TSRAM_M8
XI863 GND RBL[13] RWL[5] RWLB[5] VDD WBL[13] WBLB[13] WWLB[5] / 10TSRAM_M8
XI862 GND RBL[14] RWL[5] RWLB[5] VDD WBL[14] WBLB[14] WWLB[5] / 10TSRAM_M8
XI861 GND RBL[15] RWL[4] RWLB[4] VDD WBL[15] WBLB[15] WWLB[4] / 10TSRAM_M8
XI860 GND RBL[0] RWL[4] RWLB[4] VDD WBL[0] WBLB[0] WWLB[4] / 10TSRAM_M8
XI893 GND RBL[15] RWL[6] RWLB[6] VDD WBL[15] WBLB[15] WWLB[6] / 10TSRAM_M8
XI892 GND RBL[0] RWL[6] RWLB[6] VDD WBL[0] WBLB[0] WWLB[6] / 10TSRAM_M8
XI891 GND RBL[1] RWL[6] RWLB[6] VDD WBL[1] WBLB[1] WWLB[6] / 10TSRAM_M8
XI879 GND RBL[13] RWL[6] RWLB[6] VDD WBL[13] WBLB[13] WWLB[6] / 10TSRAM_M8
XI878 GND RBL[14] RWL[6] RWLB[6] VDD WBL[14] WBLB[14] WWLB[6] / 10TSRAM_M8
XI877 GND RBL[15] RWL[5] RWLB[5] VDD WBL[15] WBLB[15] WWLB[5] / 10TSRAM_M8
XI876 GND RBL[0] RWL[5] RWLB[5] VDD WBL[0] WBLB[0] WWLB[5] / 10TSRAM_M8
XI881 GND RBL[11] RWL[6] RWLB[6] VDD WBL[11] WBLB[11] WWLB[6] / 10TSRAM_M8
XI915 GND RBL[9] RWL[8] RWLB[8] VDD WBL[9] WBLB[9] WWLB[8] / 10TSRAM_M8
XI914 GND RBL[10] RWL[8] RWLB[8] VDD WBL[10] WBLB[10] WWLB[8] / 10TSRAM_M8
XI913 GND RBL[11] RWL[8] RWLB[8] VDD WBL[11] WBLB[11] WWLB[8] / 10TSRAM_M8
XI912 GND RBL[12] RWL[8] RWLB[8] VDD WBL[12] WBLB[12] WWLB[8] / 10TSRAM_M8
XI1027 GND RBL[9] RWL[15] RWLB[15] VDD WBL[9] WBLB[9] WWLB[15] / 10TSRAM_M8
XI1000 GND RBL[4] RWL[13] RWLB[13] VDD WBL[4] WBLB[4] WWLB[13] / 10TSRAM_M8
XI859 GND RBL[1] RWL[4] RWLB[4] VDD WBL[1] WBLB[1] WWLB[4] / 10TSRAM_M8
XI858 GND RBL[2] RWL[4] RWLB[4] VDD WBL[2] WBLB[2] WWLB[4] / 10TSRAM_M8
XI857 GND RBL[3] RWL[4] RWLB[4] VDD WBL[3] WBLB[3] WWLB[4] / 10TSRAM_M8
XI856 GND RBL[4] RWL[4] RWLB[4] VDD WBL[4] WBLB[4] WWLB[4] / 10TSRAM_M8
XI887 GND RBL[5] RWL[6] RWLB[6] VDD WBL[5] WBLB[5] WWLB[6] / 10TSRAM_M8
XI886 GND RBL[6] RWL[6] RWLB[6] VDD WBL[6] WBLB[6] WWLB[6] / 10TSRAM_M8
XI831 GND RBL[13] RWL[3] RWLB[3] VDD WBL[13] WBLB[13] WWLB[3] / 10TSRAM_M8
XI830 GND RBL[14] RWL[3] RWLB[3] VDD WBL[14] WBLB[14] WWLB[3] / 10TSRAM_M8
XI829 GND RBL[15] RWL[2] RWLB[2] VDD WBL[15] WBLB[15] WWLB[2] / 10TSRAM_M8
XI828 GND RBL[0] RWL[2] RWLB[2] VDD WBL[0] WBLB[0] WWLB[2] / 10TSRAM_M8
XI827 GND RBL[1] RWL[2] RWLB[2] VDD WBL[1] WBLB[1] WWLB[2] / 10TSRAM_M8
XI826 GND RBL[2] RWL[2] RWLB[2] VDD WBL[2] WBLB[2] WWLB[2] / 10TSRAM_M8
XI850 GND RBL[10] RWL[4] RWLB[4] VDD WBL[10] WBLB[10] WWLB[4] / 10TSRAM_M8
XI849 GND RBL[11] RWL[4] RWLB[4] VDD WBL[11] WBLB[11] WWLB[4] / 10TSRAM_M8
XI848 GND RBL[12] RWL[4] RWLB[4] VDD WBL[12] WBLB[12] WWLB[4] / 10TSRAM_M8
XI851 GND RBL[9] RWL[4] RWLB[4] VDD WBL[9] WBLB[9] WWLB[4] / 10TSRAM_M8
XI1026 GND RBL[10] RWL[15] RWLB[15] VDD WBL[10] WBLB[10] WWLB[15] / 10TSRAM_M8
XI1001 GND RBL[3] RWL[13] RWLB[13] VDD WBL[3] WBLB[3] WWLB[13] / 10TSRAM_M8
XI854 GND RBL[6] RWL[4] RWLB[4] VDD WBL[6] WBLB[6] WWLB[4] / 10TSRAM_M8
XI853 GND RBL[7] RWL[4] RWLB[4] VDD WBL[7] WBLB[7] WWLB[4] / 10TSRAM_M8
XI852 GND RBL[8] RWL[4] RWLB[4] VDD WBL[8] WBLB[8] WWLB[4] / 10TSRAM_M8
XI855 GND RBL[5] RWL[4] RWLB[4] VDD WBL[5] WBLB[5] WWLB[4] / 10TSRAM_M8
XI880 GND RBL[12] RWL[6] RWLB[6] VDD WBL[12] WBLB[12] WWLB[6] / 10TSRAM_M8
XI794 GND RBL[3] RWL[0] RWLB[0] VDD WBL[3] WBLB[3] WWLB[0] / 10TSRAM_M8
XI825 GND RBL[3] RWL[2] RWLB[2] VDD WBL[3] WBLB[3] WWLB[2] / 10TSRAM_M8
XI824 GND RBL[4] RWL[2] RWLB[2] VDD WBL[4] WBLB[4] WWLB[2] / 10TSRAM_M8
XI823 GND RBL[5] RWL[2] RWLB[2] VDD WBL[5] WBLB[5] WWLB[2] / 10TSRAM_M8
XI822 GND RBL[6] RWL[2] RWLB[2] VDD WBL[6] WBLB[6] WWLB[2] / 10TSRAM_M8
XI821 GND RBL[7] RWL[2] RWLB[2] VDD WBL[7] WBLB[7] WWLB[2] / 10TSRAM_M8
XI820 GND RBL[8] RWL[2] RWLB[2] VDD WBL[8] WBLB[8] WWLB[2] / 10TSRAM_M8
XI847 GND RBL[13] RWL[4] RWLB[4] VDD WBL[13] WBLB[13] WWLB[4] / 10TSRAM_M8
XI846 GND RBL[14] RWL[4] RWLB[4] VDD WBL[14] WBLB[14] WWLB[4] / 10TSRAM_M8
XI845 GND RBL[15] RWL[3] RWLB[3] VDD WBL[15] WBLB[15] WWLB[3] / 10TSRAM_M8
XI844 GND RBL[0] RWL[3] RWLB[3] VDD WBL[0] WBLB[0] WWLB[3] / 10TSRAM_M8
XI1025 GND RBL[11] RWL[15] RWLB[15] VDD WBL[11] WBLB[11] WWLB[15] / 10TSRAM_M8
XI1002 GND RBL[2] RWL[13] RWLB[13] VDD WBL[2] WBLB[2] WWLB[13] / 10TSRAM_M8
XI801 GND RBL[11] RWL[1] RWLB[1] VDD WBL[11] WBLB[11] WWLB[1] / 10TSRAM_M8
XI800 GND RBL[12] RWL[1] RWLB[1] VDD WBL[12] WBLB[12] WWLB[1] / 10TSRAM_M8
XI799 GND RBL[13] RWL[1] RWLB[1] VDD WBL[13] WBLB[13] WWLB[1] / 10TSRAM_M8
XI798 GND RBL[14] RWL[1] RWLB[1] VDD WBL[14] WBLB[14] WWLB[1] / 10TSRAM_M8
XI791 GND RBL[6] RWL[0] RWLB[0] VDD WBL[6] WBLB[6] WWLB[0] / 10TSRAM_M8
XI790 GND RBL[7] RWL[0] RWLB[0] VDD WBL[7] WBLB[7] WWLB[0] / 10TSRAM_M8
XI819 GND RBL[9] RWL[2] RWLB[2] VDD WBL[9] WBLB[9] WWLB[2] / 10TSRAM_M8
XI818 GND RBL[10] RWL[2] RWLB[2] VDD WBL[10] WBLB[10] WWLB[2] / 10TSRAM_M8
XI817 GND RBL[11] RWL[2] RWLB[2] VDD WBL[11] WBLB[11] WWLB[2] / 10TSRAM_M8
XI816 GND RBL[12] RWL[2] RWLB[2] VDD WBL[12] WBLB[12] WWLB[2] / 10TSRAM_M8
XI815 GND RBL[13] RWL[2] RWLB[2] VDD WBL[13] WBLB[13] WWLB[2] / 10TSRAM_M8
XI814 GND RBL[14] RWL[2] RWLB[2] VDD WBL[14] WBLB[14] WWLB[2] / 10TSRAM_M8
XI843 GND RBL[1] RWL[3] RWLB[3] VDD WBL[1] WBLB[1] WWLB[3] / 10TSRAM_M8
XI842 GND RBL[2] RWL[3] RWLB[3] VDD WBL[2] WBLB[2] WWLB[3] / 10TSRAM_M8
XI841 GND RBL[3] RWL[3] RWLB[3] VDD WBL[3] WBLB[3] WWLB[3] / 10TSRAM_M8
XI840 GND RBL[4] RWL[3] RWLB[3] VDD WBL[4] WBLB[4] WWLB[3] / 10TSRAM_M8
XI1024 GND RBL[12] RWL[15] RWLB[15] VDD WBL[12] WBLB[12] WWLB[15] / 10TSRAM_M8
XI1003 GND RBL[1] RWL[13] RWLB[13] VDD WBL[1] WBLB[1] WWLB[13] / 10TSRAM_M8
XI797 GND RBL[0] RWL[0] RWLB[0] VDD WBL[0] WBLB[0] WWLB[0] / 10TSRAM_M8
XI796 GND RBL[1] RWL[0] RWLB[0] VDD WBL[1] WBLB[1] WWLB[0] / 10TSRAM_M8
XI795 GND RBL[2] RWL[0] RWLB[0] VDD WBL[2] WBLB[2] WWLB[0] / 10TSRAM_M8
XI788 GND RBL[9] RWL[0] RWLB[0] VDD WBL[9] WBLB[9] WWLB[0] / 10TSRAM_M8
XI787 GND RBL[10] RWL[0] RWLB[0] VDD WBL[10] WBLB[10] WWLB[0] / 10TSRAM_M8
XI786 GND RBL[11] RWL[0] RWLB[0] VDD WBL[11] WBLB[11] WWLB[0] / 10TSRAM_M8
XI813 GND RBL[15] RWL[1] RWLB[1] VDD WBL[15] WBLB[15] WWLB[1] / 10TSRAM_M8
XI812 GND RBL[0] RWL[1] RWLB[1] VDD WBL[0] WBLB[0] WWLB[1] / 10TSRAM_M8
XI811 GND RBL[1] RWL[1] RWLB[1] VDD WBL[1] WBLB[1] WWLB[1] / 10TSRAM_M8
XI810 GND RBL[2] RWL[1] RWLB[1] VDD WBL[2] WBLB[2] WWLB[1] / 10TSRAM_M8
XI809 GND RBL[3] RWL[1] RWLB[1] VDD WBL[3] WBLB[3] WWLB[1] / 10TSRAM_M8
XI808 GND RBL[4] RWL[1] RWLB[1] VDD WBL[4] WBLB[4] WWLB[1] / 10TSRAM_M8
XI839 GND RBL[5] RWL[3] RWLB[3] VDD WBL[5] WBLB[5] WWLB[3] / 10TSRAM_M8
XI838 GND RBL[6] RWL[3] RWLB[3] VDD WBL[6] WBLB[6] WWLB[3] / 10TSRAM_M8
XI837 GND RBL[7] RWL[3] RWLB[3] VDD WBL[7] WBLB[7] WWLB[3] / 10TSRAM_M8
XI836 GND RBL[8] RWL[3] RWLB[3] VDD WBL[8] WBLB[8] WWLB[3] / 10TSRAM_M8
XI1023 GND RBL[13] RWL[15] RWLB[15] VDD WBL[13] WBLB[13] WWLB[15] / 10TSRAM_M8
XI1004 GND RBL[0] RWL[13] RWLB[13] VDD WBL[0] WBLB[0] WWLB[13] / 10TSRAM_M8
XI793 GND RBL[4] RWL[0] RWLB[0] VDD WBL[4] WBLB[4] WWLB[0] / 10TSRAM_M8
XI792 GND RBL[5] RWL[0] RWLB[0] VDD WBL[5] WBLB[5] WWLB[0] / 10TSRAM_M8
XI784 GND RBL[13] RWL[0] RWLB[0] VDD WBL[13] WBLB[13] WWLB[0] / 10TSRAM_M8
XI783 GND RBL[14] RWL[0] RWLB[0] VDD WBL[14] WBLB[14] WWLB[0] / 10TSRAM_M8
XI782 GND RBL[15] RWL[0] RWLB[0] VDD WBL[15] WBLB[15] WWLB[0] / 10TSRAM_M8
XI785 GND RBL[12] RWL[0] RWLB[0] VDD WBL[12] WBLB[12] WWLB[0] / 10TSRAM_M8
XI806 GND RBL[6] RWL[1] RWLB[1] VDD WBL[6] WBLB[6] WWLB[1] / 10TSRAM_M8
XI805 GND RBL[7] RWL[1] RWLB[1] VDD WBL[7] WBLB[7] WWLB[1] / 10TSRAM_M8
XI804 GND RBL[8] RWL[1] RWLB[1] VDD WBL[8] WBLB[8] WWLB[1] / 10TSRAM_M8
XI803 GND RBL[9] RWL[1] RWLB[1] VDD WBL[9] WBLB[9] WWLB[1] / 10TSRAM_M8
XI802 GND RBL[10] RWL[1] RWLB[1] VDD WBL[10] WBLB[10] WWLB[1] / 10TSRAM_M8
XI807 GND RBL[5] RWL[1] RWLB[1] VDD WBL[5] WBLB[5] WWLB[1] / 10TSRAM_M8
XI835 GND RBL[9] RWL[3] RWLB[3] VDD WBL[9] WBLB[9] WWLB[3] / 10TSRAM_M8
XI834 GND RBL[10] RWL[3] RWLB[3] VDD WBL[10] WBLB[10] WWLB[3] / 10TSRAM_M8
XI833 GND RBL[11] RWL[3] RWLB[3] VDD WBL[11] WBLB[11] WWLB[3] / 10TSRAM_M8
XI832 GND RBL[12] RWL[3] RWLB[3] VDD WBL[12] WBLB[12] WWLB[3] / 10TSRAM_M8
XI1022 GND RBL[14] RWL[15] RWLB[15] VDD WBL[14] WBLB[14] WWLB[15] / 10TSRAM_M8
XI1005 GND RBL[15] RWL[13] RWLB[13] VDD WBL[15] WBLB[15] WWLB[13] / 10TSRAM_M8
XI789 GND RBL[8] RWL[0] RWLB[0] VDD WBL[8] WBLB[8] WWLB[0] / 10TSRAM_M8
.ENDS

