* File: /home/wjin/dmtalen/sram/10TSRAM_PEX/16x16_10T_new.pex.netlist
* Created: Mon Aug 14 10:51:10 2017
* Program "Calibre xRC"
* Version "v2011.3_18.12"
* 
.include "/home/wjin/dmtalen/sram/10TSRAM_PEX/16x16_10T_new.pex.netlist.pex"
.subckt array16x16_10T_new  wwlb<15> wwlb<14> wwlb<13> wwlb<12> wwlb<11> wwlb<10>
+ wwlb<9> wwlb<8> wwlb<7> wwlb<6> wwlb<5> wwlb<4> wwlb<3> wwlb<2> wwlb<1>
+ wwlb<0> rwl<15> rwl<14> rwl<13> rwl<12> rwl<11> rwl<10> rwl<9> rwl<8> rwl<7>
+ rwl<6> rwl<5> rwl<4> rwl<3> rwl<2> rwl<1> rwl<0> rwlb<15> rwlb<14> rwlb<13>
+ rwlb<12> rwlb<11> rwlb<10> rwlb<9> rwlb<8> rwlb<7> rwlb<6> rwlb<5> rwlb<4>
+ rwlb<3> rwlb<2> rwlb<1> rwlb<0> wbl<15> wbl<14> wbl<13> wbl<12> wbl<11>
+ wbl<10> wbl<9> wbl<8> wbl<7> wbl<6> wbl<5> wbl<4> wbl<3> wbl<2> wbl<1> wbl<0> + wblb<15> wblb<14> wblb<13> wblb<12> wblb<11> wblb<10> wblb<9> wblb<8> wblb<7>
+ wblb<6> wblb<5> wblb<4> wblb<3> wblb<2> wblb<1> wblb<0> rbl<15> rbl<14>
+ rbl<13> rbl<12> rbl<11> rbl<10> rbl<9> rbl<8> rbl<7> rbl<6> rbl<5> rbl<4>
+ rbl<3> rbl<2> rbl<1> rbl<0>
* 
* WBLB<0>	WBLB<0>
* WBL<0>	WBL<0>
* WBL<1>	WBL<1>
* WBLB<1>	WBLB<1>
* WBLB<2>	WBLB<2>
* WBL<2>	WBL<2>
* WBL<3>	WBL<3>
* WBLB<3>	WBLB<3>
* WBLB<4>	WBLB<4>
* WBL<4>	WBL<4>
* WBL<5>	WBL<5>
* WBLB<5>	WBLB<5>
* WBLB<6>	WBLB<6>
* WBL<6>	WBL<6>
* WBL<7>	WBL<7>
* WBLB<7>	WBLB<7>
* WBLB<8>	WBLB<8>
* WBL<8>	WBL<8>
* WBL<9>	WBL<9>
* WBLB<9>	WBLB<9>
* WBLB<10>	WBLB<10>
* WBL<10>	WBL<10>
* WBL<11>	WBL<11>
* WBLB<11>	WBLB<11>
* WBLB<12>	WBLB<12>
* WBL<12>	WBL<12>
* WBL<13>	WBL<13>
* WBLB<13>	WBLB<13>
* WBLB<14>	WBLB<14>
* WBL<14>	WBL<14>
* WBL<15>	WBL<15>
* WBLB<15>	WBLB<15>
* RWL<7>	RWL<7>
* RWL<6>	RWL<6>
* RWL<5>	RWL<5>
* RWL<4>	RWL<4>
* RWL<3>	RWL<3>
* RWL<2>	RWL<2>
* RWL<1>	RWL<1>
* RWL<0>	RWL<0>
* WWLB<7>	WWLB<7>
* WWLB<6>	WWLB<6>
* WWLB<5>	WWLB<5>
* WWLB<4>	WWLB<4>
* WWLB<3>	WWLB<3>
* WWLB<2>	WWLB<2>
* WWLB<1>	WWLB<1>
* WWLB<0>	WWLB<0>
* RWL<15>	RWL<15>
* RWL<14>	RWL<14>
* RWL<13>	RWL<13>
* RWL<12>	RWL<12>
* RWL<11>	RWL<11>
* RWL<10>	RWL<10>
* RWL<9>	RWL<9>
* RWL<8>	RWL<8>
* WWLB<15>	WWLB<15>
* WWLB<14>	WWLB<14>
* WWLB<13>	WWLB<13>
* WWLB<12>	WWLB<12>
* WWLB<11>	WWLB<11>
* WWLB<10>	WWLB<10>
* WWLB<9>	WWLB<9>
* WWLB<8>	WWLB<8>
* GND	GND
* RWLB<7>	RWLB<7>
* RWLB<6>	RWLB<6>
* RWLB<5>	RWLB<5>
* RWLB<4>	RWLB<4>
* RWLB<3>	RWLB<3>
* RWLB<2>	RWLB<2>
* RWLB<1>	RWLB<1>
* RWLB<0>	RWLB<0>
* RWLB<15>	RWLB<15>
* RWLB<14>	RWLB<14>
* RWLB<13>	RWLB<13>
* RWLB<12>	RWLB<12>
* RWLB<11>	RWLB<11>
* RWLB<10>	RWLB<10>
* RWLB<9>	RWLB<9>
* RWLB<8>	RWLB<8>
* VDD	VDD
* RBL<0>	RBL<0>
* RBL<1>	RBL<1>
* RBL<2>	RBL<2>
* RBL<3>	RBL<3>
* RBL<4>	RBL<4>
* RBL<5>	RBL<5>
* RBL<6>	RBL<6>
* RBL<7>	RBL<7>
* RBL<8>	RBL<8>
* RBL<9>	RBL<9>
* RBL<10>	RBL<10>
* RBL<11>	RBL<11>
* RBL<12>	RBL<12>
* RBL<13>	RBL<13>
* RBL<14>	RBL<14>
* RBL<15>	RBL<15>
mXI1006/MM8 N_XI1006/NET08_XI1006/MM8_d N_RWL<14>_XI1006/MM8_g
+ N_RBL<14>_XI1006/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1006/MM7 N_XI1006/NET08_XI1006/MM7_d N_XI1006/QB_XI1006/MM7_g
+ N_GND_XI1006/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1006/MM10 N_WBL<14>_XI1006/MM10_d N_WWLB<14>_XI1006/MM10_g
+ N_XI1006/Q_XI1006/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1006/MM11 N_WBLB<14>_XI1006/MM11_d N_WWLB<14>_XI1006/MM11_g
+ N_XI1006/QB_XI1006/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1006/MM1 N_XI1006/Q_XI1006/MM1_d N_XI1006/QB_XI1006/MM1_g N_GND_XI1006/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1006/MM0 N_XI1006/QB_XI1006/MM0_d N_XI1006/Q_XI1006/MM0_g N_GND_XI1006/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1006/MM9 N_XI1006/NET08_XI1006/MM9_d N_RWLB<14>_XI1006/MM9_g
+ N_RBL<14>_XI1006/MM9_s N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1006/MM6 N_XI1006/NET08_XI1006/MM6_d N_XI1006/QB_XI1006/MM6_g
+ N_VDD_XI1006/MM6_s N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1006/MM5 N_XI1006/Q_XI1006/MM5_d N_XI1006/QB_XI1006/MM5_g N_VDD_XI1006/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1006/MM4 N_XI1006/QB_XI1006/MM4_d N_XI1006/Q_XI1006/MM4_g N_VDD_XI1006/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1020/MM8 N_XI1020/NET08_XI1020/MM8_d N_RWL<14>_XI1020/MM8_g
+ N_RBL<0>_XI1020/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1020/MM7 N_XI1020/NET08_XI1020/MM7_d N_XI1020/QB_XI1020/MM7_g
+ N_GND_XI1020/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1020/MM10 N_WBL<0>_XI1020/MM10_d N_WWLB<14>_XI1020/MM10_g
+ N_XI1020/Q_XI1020/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1020/MM11 N_WBLB<0>_XI1020/MM11_d N_WWLB<14>_XI1020/MM11_g
+ N_XI1020/QB_XI1020/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1020/MM1 N_XI1020/Q_XI1020/MM1_d N_XI1020/QB_XI1020/MM1_g N_GND_XI1020/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1020/MM0 N_XI1020/QB_XI1020/MM0_d N_XI1020/Q_XI1020/MM0_g N_GND_XI1020/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1020/MM9 N_XI1020/NET08_XI1020/MM9_d N_RWLB<14>_XI1020/MM9_g
+ N_RBL<0>_XI1020/MM9_s N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1020/MM6 N_XI1020/NET08_XI1020/MM6_d N_XI1020/QB_XI1020/MM6_g
+ N_VDD_XI1020/MM6_s N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1020/MM5 N_XI1020/Q_XI1020/MM5_d N_XI1020/QB_XI1020/MM5_g N_VDD_XI1020/MM5_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1020/MM4 N_XI1020/QB_XI1020/MM4_d N_XI1020/Q_XI1020/MM4_g N_VDD_XI1020/MM4_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1019/MM8 N_XI1019/NET08_XI1019/MM8_d N_RWL<14>_XI1019/MM8_g
+ N_RBL<1>_XI1019/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1019/MM7 N_XI1019/NET08_XI1019/MM7_d N_XI1019/QB_XI1019/MM7_g
+ N_GND_XI1019/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1019/MM10 N_WBL<1>_XI1019/MM10_d N_WWLB<14>_XI1019/MM10_g
+ N_XI1019/Q_XI1019/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1019/MM11 N_WBLB<1>_XI1019/MM11_d N_WWLB<14>_XI1019/MM11_g
+ N_XI1019/QB_XI1019/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1019/MM1 N_XI1019/Q_XI1019/MM1_d N_XI1019/QB_XI1019/MM1_g N_GND_XI1019/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1019/MM0 N_XI1019/QB_XI1019/MM0_d N_XI1019/Q_XI1019/MM0_g N_GND_XI1019/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1019/MM9 N_XI1019/NET08_XI1019/MM9_d N_RWLB<14>_XI1019/MM9_g
+ N_RBL<1>_XI1019/MM9_s N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1019/MM6 N_XI1019/NET08_XI1019/MM6_d N_XI1019/QB_XI1019/MM6_g
+ N_VDD_XI1019/MM6_s N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1019/MM5 N_XI1019/Q_XI1019/MM5_d N_XI1019/QB_XI1019/MM5_g N_VDD_XI1019/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1019/MM4 N_XI1019/QB_XI1019/MM4_d N_XI1019/Q_XI1019/MM4_g N_VDD_XI1019/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1018/MM8 N_XI1018/NET08_XI1018/MM8_d N_RWL<14>_XI1018/MM8_g
+ N_RBL<2>_XI1018/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1018/MM7 N_XI1018/NET08_XI1018/MM7_d N_XI1018/QB_XI1018/MM7_g
+ N_GND_XI1018/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1018/MM10 N_WBL<2>_XI1018/MM10_d N_WWLB<14>_XI1018/MM10_g
+ N_XI1018/Q_XI1018/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1018/MM11 N_WBLB<2>_XI1018/MM11_d N_WWLB<14>_XI1018/MM11_g
+ N_XI1018/QB_XI1018/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1018/MM1 N_XI1018/Q_XI1018/MM1_d N_XI1018/QB_XI1018/MM1_g N_GND_XI1018/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1018/MM0 N_XI1018/QB_XI1018/MM0_d N_XI1018/Q_XI1018/MM0_g N_GND_XI1018/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1018/MM9 N_XI1018/NET08_XI1018/MM9_d N_RWLB<14>_XI1018/MM9_g
+ N_RBL<2>_XI1018/MM9_s N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1018/MM6 N_XI1018/NET08_XI1018/MM6_d N_XI1018/QB_XI1018/MM6_g
+ N_VDD_XI1018/MM6_s N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1018/MM5 N_XI1018/Q_XI1018/MM5_d N_XI1018/QB_XI1018/MM5_g N_VDD_XI1018/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1018/MM4 N_XI1018/QB_XI1018/MM4_d N_XI1018/Q_XI1018/MM4_g N_VDD_XI1018/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1017/MM8 N_XI1017/NET08_XI1017/MM8_d N_RWL<14>_XI1017/MM8_g
+ N_RBL<3>_XI1017/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1017/MM7 N_XI1017/NET08_XI1017/MM7_d N_XI1017/QB_XI1017/MM7_g
+ N_GND_XI1017/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1017/MM10 N_WBL<3>_XI1017/MM10_d N_WWLB<14>_XI1017/MM10_g
+ N_XI1017/Q_XI1017/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1017/MM11 N_WBLB<3>_XI1017/MM11_d N_WWLB<14>_XI1017/MM11_g
+ N_XI1017/QB_XI1017/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1017/MM1 N_XI1017/Q_XI1017/MM1_d N_XI1017/QB_XI1017/MM1_g N_GND_XI1017/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1017/MM0 N_XI1017/QB_XI1017/MM0_d N_XI1017/Q_XI1017/MM0_g N_GND_XI1017/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1017/MM9 N_XI1017/NET08_XI1017/MM9_d N_RWLB<14>_XI1017/MM9_g
+ N_RBL<3>_XI1017/MM9_s N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1017/MM6 N_XI1017/NET08_XI1017/MM6_d N_XI1017/QB_XI1017/MM6_g
+ N_VDD_XI1017/MM6_s N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1017/MM5 N_XI1017/Q_XI1017/MM5_d N_XI1017/QB_XI1017/MM5_g N_VDD_XI1017/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1017/MM4 N_XI1017/QB_XI1017/MM4_d N_XI1017/Q_XI1017/MM4_g N_VDD_XI1017/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1016/MM8 N_XI1016/NET08_XI1016/MM8_d N_RWL<14>_XI1016/MM8_g
+ N_RBL<4>_XI1016/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1016/MM7 N_XI1016/NET08_XI1016/MM7_d N_XI1016/QB_XI1016/MM7_g
+ N_GND_XI1016/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1016/MM10 N_WBL<4>_XI1016/MM10_d N_WWLB<14>_XI1016/MM10_g
+ N_XI1016/Q_XI1016/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1016/MM11 N_WBLB<4>_XI1016/MM11_d N_WWLB<14>_XI1016/MM11_g
+ N_XI1016/QB_XI1016/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1016/MM1 N_XI1016/Q_XI1016/MM1_d N_XI1016/QB_XI1016/MM1_g N_GND_XI1016/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1016/MM0 N_XI1016/QB_XI1016/MM0_d N_XI1016/Q_XI1016/MM0_g N_GND_XI1016/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1016/MM9 N_XI1016/NET08_XI1016/MM9_d N_RWLB<14>_XI1016/MM9_g
+ N_RBL<4>_XI1016/MM9_s N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1016/MM6 N_XI1016/NET08_XI1016/MM6_d N_XI1016/QB_XI1016/MM6_g
+ N_VDD_XI1016/MM6_s N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1016/MM5 N_XI1016/Q_XI1016/MM5_d N_XI1016/QB_XI1016/MM5_g N_VDD_XI1016/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1016/MM4 N_XI1016/QB_XI1016/MM4_d N_XI1016/Q_XI1016/MM4_g N_VDD_XI1016/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1015/MM8 N_XI1015/NET08_XI1015/MM8_d N_RWL<14>_XI1015/MM8_g
+ N_RBL<5>_XI1015/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1015/MM7 N_XI1015/NET08_XI1015/MM7_d N_XI1015/QB_XI1015/MM7_g
+ N_GND_XI1015/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1015/MM10 N_WBL<5>_XI1015/MM10_d N_WWLB<14>_XI1015/MM10_g
+ N_XI1015/Q_XI1015/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1015/MM11 N_WBLB<5>_XI1015/MM11_d N_WWLB<14>_XI1015/MM11_g
+ N_XI1015/QB_XI1015/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1015/MM1 N_XI1015/Q_XI1015/MM1_d N_XI1015/QB_XI1015/MM1_g N_GND_XI1015/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1015/MM0 N_XI1015/QB_XI1015/MM0_d N_XI1015/Q_XI1015/MM0_g N_GND_XI1015/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1015/MM9 N_XI1015/NET08_XI1015/MM9_d N_RWLB<14>_XI1015/MM9_g
+ N_RBL<5>_XI1015/MM9_s N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1015/MM6 N_XI1015/NET08_XI1015/MM6_d N_XI1015/QB_XI1015/MM6_g
+ N_VDD_XI1015/MM6_s N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1015/MM5 N_XI1015/Q_XI1015/MM5_d N_XI1015/QB_XI1015/MM5_g N_VDD_XI1015/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1015/MM4 N_XI1015/QB_XI1015/MM4_d N_XI1015/Q_XI1015/MM4_g N_VDD_XI1015/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1014/MM8 N_XI1014/NET08_XI1014/MM8_d N_RWL<14>_XI1014/MM8_g
+ N_RBL<6>_XI1014/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1014/MM7 N_XI1014/NET08_XI1014/MM7_d N_XI1014/QB_XI1014/MM7_g
+ N_GND_XI1014/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1014/MM10 N_WBL<6>_XI1014/MM10_d N_WWLB<14>_XI1014/MM10_g
+ N_XI1014/Q_XI1014/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1014/MM11 N_WBLB<6>_XI1014/MM11_d N_WWLB<14>_XI1014/MM11_g
+ N_XI1014/QB_XI1014/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1014/MM1 N_XI1014/Q_XI1014/MM1_d N_XI1014/QB_XI1014/MM1_g N_GND_XI1014/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1014/MM0 N_XI1014/QB_XI1014/MM0_d N_XI1014/Q_XI1014/MM0_g N_GND_XI1014/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1014/MM9 N_XI1014/NET08_XI1014/MM9_d N_RWLB<14>_XI1014/MM9_g
+ N_RBL<6>_XI1014/MM9_s N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1014/MM6 N_XI1014/NET08_XI1014/MM6_d N_XI1014/QB_XI1014/MM6_g
+ N_VDD_XI1014/MM6_s N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1014/MM5 N_XI1014/Q_XI1014/MM5_d N_XI1014/QB_XI1014/MM5_g N_VDD_XI1014/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1014/MM4 N_XI1014/QB_XI1014/MM4_d N_XI1014/Q_XI1014/MM4_g N_VDD_XI1014/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1013/MM8 N_XI1013/NET08_XI1013/MM8_d N_RWL<14>_XI1013/MM8_g
+ N_RBL<7>_XI1013/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1013/MM7 N_XI1013/NET08_XI1013/MM7_d N_XI1013/QB_XI1013/MM7_g
+ N_GND_XI1013/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1013/MM10 N_WBL<7>_XI1013/MM10_d N_WWLB<14>_XI1013/MM10_g
+ N_XI1013/Q_XI1013/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1013/MM11 N_WBLB<7>_XI1013/MM11_d N_WWLB<14>_XI1013/MM11_g
+ N_XI1013/QB_XI1013/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1013/MM1 N_XI1013/Q_XI1013/MM1_d N_XI1013/QB_XI1013/MM1_g N_GND_XI1013/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1013/MM0 N_XI1013/QB_XI1013/MM0_d N_XI1013/Q_XI1013/MM0_g N_GND_XI1013/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1013/MM9 N_XI1013/NET08_XI1013/MM9_d N_RWLB<14>_XI1013/MM9_g
+ N_RBL<7>_XI1013/MM9_s N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1013/MM6 N_XI1013/NET08_XI1013/MM6_d N_XI1013/QB_XI1013/MM6_g
+ N_VDD_XI1013/MM6_s N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1013/MM5 N_XI1013/Q_XI1013/MM5_d N_XI1013/QB_XI1013/MM5_g N_VDD_XI1013/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1013/MM4 N_XI1013/QB_XI1013/MM4_d N_XI1013/Q_XI1013/MM4_g N_VDD_XI1013/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1012/MM8 N_XI1012/NET08_XI1012/MM8_d N_RWL<14>_XI1012/MM8_g
+ N_RBL<8>_XI1012/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1012/MM7 N_XI1012/NET08_XI1012/MM7_d N_XI1012/QB_XI1012/MM7_g
+ N_GND_XI1012/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1012/MM10 N_WBL<8>_XI1012/MM10_d N_WWLB<14>_XI1012/MM10_g
+ N_XI1012/Q_XI1012/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1012/MM11 N_WBLB<8>_XI1012/MM11_d N_WWLB<14>_XI1012/MM11_g
+ N_XI1012/QB_XI1012/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1012/MM1 N_XI1012/Q_XI1012/MM1_d N_XI1012/QB_XI1012/MM1_g N_GND_XI1012/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1012/MM0 N_XI1012/QB_XI1012/MM0_d N_XI1012/Q_XI1012/MM0_g N_GND_XI1012/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1012/MM9 N_XI1012/NET08_XI1012/MM9_d N_RWLB<14>_XI1012/MM9_g
+ N_RBL<8>_XI1012/MM9_s N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1012/MM6 N_XI1012/NET08_XI1012/MM6_d N_XI1012/QB_XI1012/MM6_g
+ N_VDD_XI1012/MM6_s N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1012/MM5 N_XI1012/Q_XI1012/MM5_d N_XI1012/QB_XI1012/MM5_g N_VDD_XI1012/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1012/MM4 N_XI1012/QB_XI1012/MM4_d N_XI1012/Q_XI1012/MM4_g N_VDD_XI1012/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1011/MM8 N_XI1011/NET08_XI1011/MM8_d N_RWL<14>_XI1011/MM8_g
+ N_RBL<9>_XI1011/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1011/MM7 N_XI1011/NET08_XI1011/MM7_d N_XI1011/QB_XI1011/MM7_g
+ N_GND_XI1011/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1011/MM10 N_WBL<9>_XI1011/MM10_d N_WWLB<14>_XI1011/MM10_g
+ N_XI1011/Q_XI1011/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1011/MM11 N_WBLB<9>_XI1011/MM11_d N_WWLB<14>_XI1011/MM11_g
+ N_XI1011/QB_XI1011/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1011/MM1 N_XI1011/Q_XI1011/MM1_d N_XI1011/QB_XI1011/MM1_g N_GND_XI1011/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1011/MM0 N_XI1011/QB_XI1011/MM0_d N_XI1011/Q_XI1011/MM0_g N_GND_XI1011/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1011/MM9 N_XI1011/NET08_XI1011/MM9_d N_RWLB<14>_XI1011/MM9_g
+ N_RBL<9>_XI1011/MM9_s N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1011/MM6 N_XI1011/NET08_XI1011/MM6_d N_XI1011/QB_XI1011/MM6_g
+ N_VDD_XI1011/MM6_s N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1011/MM5 N_XI1011/Q_XI1011/MM5_d N_XI1011/QB_XI1011/MM5_g N_VDD_XI1011/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1011/MM4 N_XI1011/QB_XI1011/MM4_d N_XI1011/Q_XI1011/MM4_g N_VDD_XI1011/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1010/MM8 N_XI1010/NET08_XI1010/MM8_d N_RWL<14>_XI1010/MM8_g
+ N_RBL<10>_XI1010/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1010/MM7 N_XI1010/NET08_XI1010/MM7_d N_XI1010/QB_XI1010/MM7_g
+ N_GND_XI1010/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1010/MM10 N_WBL<10>_XI1010/MM10_d N_WWLB<14>_XI1010/MM10_g
+ N_XI1010/Q_XI1010/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1010/MM11 N_WBLB<10>_XI1010/MM11_d N_WWLB<14>_XI1010/MM11_g
+ N_XI1010/QB_XI1010/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1010/MM1 N_XI1010/Q_XI1010/MM1_d N_XI1010/QB_XI1010/MM1_g N_GND_XI1010/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1010/MM0 N_XI1010/QB_XI1010/MM0_d N_XI1010/Q_XI1010/MM0_g N_GND_XI1010/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1010/MM9 N_XI1010/NET08_XI1010/MM9_d N_RWLB<14>_XI1010/MM9_g
+ N_RBL<10>_XI1010/MM9_s N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1010/MM6 N_XI1010/NET08_XI1010/MM6_d N_XI1010/QB_XI1010/MM6_g
+ N_VDD_XI1010/MM6_s N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1010/MM5 N_XI1010/Q_XI1010/MM5_d N_XI1010/QB_XI1010/MM5_g N_VDD_XI1010/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1010/MM4 N_XI1010/QB_XI1010/MM4_d N_XI1010/Q_XI1010/MM4_g N_VDD_XI1010/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1009/MM8 N_XI1009/NET08_XI1009/MM8_d N_RWL<14>_XI1009/MM8_g
+ N_RBL<11>_XI1009/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1009/MM7 N_XI1009/NET08_XI1009/MM7_d N_XI1009/QB_XI1009/MM7_g
+ N_GND_XI1009/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1009/MM10 N_WBL<11>_XI1009/MM10_d N_WWLB<14>_XI1009/MM10_g
+ N_XI1009/Q_XI1009/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1009/MM11 N_WBLB<11>_XI1009/MM11_d N_WWLB<14>_XI1009/MM11_g
+ N_XI1009/QB_XI1009/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1009/MM1 N_XI1009/Q_XI1009/MM1_d N_XI1009/QB_XI1009/MM1_g N_GND_XI1009/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1009/MM0 N_XI1009/QB_XI1009/MM0_d N_XI1009/Q_XI1009/MM0_g N_GND_XI1009/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1009/MM9 N_XI1009/NET08_XI1009/MM9_d N_RWLB<14>_XI1009/MM9_g
+ N_RBL<11>_XI1009/MM9_s N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1009/MM6 N_XI1009/NET08_XI1009/MM6_d N_XI1009/QB_XI1009/MM6_g
+ N_VDD_XI1009/MM6_s N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1009/MM5 N_XI1009/Q_XI1009/MM5_d N_XI1009/QB_XI1009/MM5_g N_VDD_XI1009/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1009/MM4 N_XI1009/QB_XI1009/MM4_d N_XI1009/Q_XI1009/MM4_g N_VDD_XI1009/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1008/MM8 N_XI1008/NET08_XI1008/MM8_d N_RWL<14>_XI1008/MM8_g
+ N_RBL<12>_XI1008/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1008/MM7 N_XI1008/NET08_XI1008/MM7_d N_XI1008/QB_XI1008/MM7_g
+ N_GND_XI1008/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1008/MM10 N_WBL<12>_XI1008/MM10_d N_WWLB<14>_XI1008/MM10_g
+ N_XI1008/Q_XI1008/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1008/MM11 N_WBLB<12>_XI1008/MM11_d N_WWLB<14>_XI1008/MM11_g
+ N_XI1008/QB_XI1008/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1008/MM1 N_XI1008/Q_XI1008/MM1_d N_XI1008/QB_XI1008/MM1_g N_GND_XI1008/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1008/MM0 N_XI1008/QB_XI1008/MM0_d N_XI1008/Q_XI1008/MM0_g N_GND_XI1008/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1008/MM9 N_XI1008/NET08_XI1008/MM9_d N_RWLB<14>_XI1008/MM9_g
+ N_RBL<12>_XI1008/MM9_s N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1008/MM6 N_XI1008/NET08_XI1008/MM6_d N_XI1008/QB_XI1008/MM6_g
+ N_VDD_XI1008/MM6_s N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1008/MM5 N_XI1008/Q_XI1008/MM5_d N_XI1008/QB_XI1008/MM5_g N_VDD_XI1008/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1008/MM4 N_XI1008/QB_XI1008/MM4_d N_XI1008/Q_XI1008/MM4_g N_VDD_XI1008/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1007/MM8 N_XI1007/NET08_XI1007/MM8_d N_RWL<14>_XI1007/MM8_g
+ N_RBL<13>_XI1007/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1007/MM7 N_XI1007/NET08_XI1007/MM7_d N_XI1007/QB_XI1007/MM7_g
+ N_GND_XI1007/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1007/MM10 N_WBL<13>_XI1007/MM10_d N_WWLB<14>_XI1007/MM10_g
+ N_XI1007/Q_XI1007/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1007/MM11 N_WBLB<13>_XI1007/MM11_d N_WWLB<14>_XI1007/MM11_g
+ N_XI1007/QB_XI1007/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1007/MM1 N_XI1007/Q_XI1007/MM1_d N_XI1007/QB_XI1007/MM1_g N_GND_XI1007/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1007/MM0 N_XI1007/QB_XI1007/MM0_d N_XI1007/Q_XI1007/MM0_g N_GND_XI1007/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1007/MM9 N_XI1007/NET08_XI1007/MM9_d N_RWLB<14>_XI1007/MM9_g
+ N_RBL<13>_XI1007/MM9_s N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1007/MM6 N_XI1007/NET08_XI1007/MM6_d N_XI1007/QB_XI1007/MM6_g
+ N_VDD_XI1007/MM6_s N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1007/MM5 N_XI1007/Q_XI1007/MM5_d N_XI1007/QB_XI1007/MM5_g N_VDD_XI1007/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1007/MM4 N_XI1007/QB_XI1007/MM4_d N_XI1007/Q_XI1007/MM4_g N_VDD_XI1007/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1021/MM8 N_XI1021/NET08_XI1021/MM8_d N_RWL<14>_XI1021/MM8_g
+ N_RBL<15>_XI1021/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1021/MM7 N_XI1021/NET08_XI1021/MM7_d N_XI1021/QB_XI1021/MM7_g
+ N_GND_XI1021/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1021/MM10 N_WBL<15>_XI1021/MM10_d N_WWLB<14>_XI1021/MM10_g
+ N_XI1021/Q_XI1021/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1021/MM11 N_WBLB<15>_XI1021/MM11_d N_WWLB<14>_XI1021/MM11_g
+ N_XI1021/QB_XI1021/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1021/MM1 N_XI1021/Q_XI1021/MM1_d N_XI1021/QB_XI1021/MM1_g N_GND_XI1021/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1021/MM0 N_XI1021/QB_XI1021/MM0_d N_XI1021/Q_XI1021/MM0_g N_GND_XI1021/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1021/MM9 N_XI1021/NET08_XI1021/MM9_d N_RWLB<14>_XI1021/MM9_g
+ N_RBL<15>_XI1021/MM9_s N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1021/MM6 N_XI1021/NET08_XI1021/MM6_d N_XI1021/QB_XI1021/MM6_g
+ N_VDD_XI1021/MM6_s N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1021/MM5 N_XI1021/Q_XI1021/MM5_d N_XI1021/QB_XI1021/MM5_g N_VDD_XI1021/MM5_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1021/MM4 N_XI1021/QB_XI1021/MM4_d N_XI1021/Q_XI1021/MM4_g N_VDD_XI1021/MM4_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1037/MM8 N_XI1037/NET08_XI1037/MM8_d N_RWL<15>_XI1037/MM8_g
+ N_RBL<15>_XI1037/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1037/MM7 N_XI1037/NET08_XI1037/MM7_d N_XI1037/QB_XI1037/MM7_g
+ N_GND_XI1037/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1037/MM10 N_WBL<15>_XI1037/MM10_d N_WWLB<15>_XI1037/MM10_g
+ N_XI1037/Q_XI1037/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1037/MM11 N_WBLB<15>_XI1037/MM11_d N_WWLB<15>_XI1037/MM11_g
+ N_XI1037/QB_XI1037/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1037/MM1 N_XI1037/Q_XI1037/MM1_d N_XI1037/QB_XI1037/MM1_g N_GND_XI1037/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1037/MM0 N_XI1037/QB_XI1037/MM0_d N_XI1037/Q_XI1037/MM0_g N_GND_XI1037/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1037/MM9 N_XI1037/NET08_XI1037/MM9_d N_RWLB<15>_XI1037/MM9_g
+ N_RBL<15>_XI1037/MM9_s N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1037/MM6 N_XI1037/NET08_XI1037/MM6_d N_XI1037/QB_XI1037/MM6_g
+ N_VDD_XI1037/MM6_s N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1037/MM5 N_XI1037/Q_XI1037/MM5_d N_XI1037/QB_XI1037/MM5_g N_VDD_XI1037/MM5_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1037/MM4 N_XI1037/QB_XI1037/MM4_d N_XI1037/Q_XI1037/MM4_g N_VDD_XI1037/MM4_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1036/MM8 N_XI1036/NET08_XI1036/MM8_d N_RWL<15>_XI1036/MM8_g
+ N_RBL<0>_XI1036/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1036/MM7 N_XI1036/NET08_XI1036/MM7_d N_XI1036/QB_XI1036/MM7_g
+ N_GND_XI1036/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1036/MM10 N_WBL<0>_XI1036/MM10_d N_WWLB<15>_XI1036/MM10_g
+ N_XI1036/Q_XI1036/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1036/MM11 N_WBLB<0>_XI1036/MM11_d N_WWLB<15>_XI1036/MM11_g
+ N_XI1036/QB_XI1036/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1036/MM1 N_XI1036/Q_XI1036/MM1_d N_XI1036/QB_XI1036/MM1_g N_GND_XI1036/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1036/MM0 N_XI1036/QB_XI1036/MM0_d N_XI1036/Q_XI1036/MM0_g N_GND_XI1036/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1036/MM9 N_XI1036/NET08_XI1036/MM9_d N_RWLB<15>_XI1036/MM9_g
+ N_RBL<0>_XI1036/MM9_s N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1036/MM6 N_XI1036/NET08_XI1036/MM6_d N_XI1036/QB_XI1036/MM6_g
+ N_VDD_XI1036/MM6_s N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1036/MM5 N_XI1036/Q_XI1036/MM5_d N_XI1036/QB_XI1036/MM5_g N_VDD_XI1036/MM5_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1036/MM4 N_XI1036/QB_XI1036/MM4_d N_XI1036/Q_XI1036/MM4_g N_VDD_XI1036/MM4_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI984/MM8 N_XI984/NET08_XI984/MM8_d N_RWL<12>_XI984/MM8_g N_RBL<4>_XI984/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI984/MM7 N_XI984/NET08_XI984/MM7_d N_XI984/QB_XI984/MM7_g N_GND_XI984/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI984/MM10 N_WBL<4>_XI984/MM10_d N_WWLB<12>_XI984/MM10_g N_XI984/Q_XI984/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI984/MM11 N_WBLB<4>_XI984/MM11_d N_WWLB<12>_XI984/MM11_g
+ N_XI984/QB_XI984/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI984/MM1 N_XI984/Q_XI984/MM1_d N_XI984/QB_XI984/MM1_g N_GND_XI984/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI984/MM0 N_XI984/QB_XI984/MM0_d N_XI984/Q_XI984/MM0_g N_GND_XI984/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI984/MM9 N_XI984/NET08_XI984/MM9_d N_RWLB<12>_XI984/MM9_g N_RBL<4>_XI984/MM9_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI984/MM6 N_XI984/NET08_XI984/MM6_d N_XI984/QB_XI984/MM6_g N_VDD_XI984/MM6_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI984/MM5 N_XI984/Q_XI984/MM5_d N_XI984/QB_XI984/MM5_g N_VDD_XI984/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI984/MM4 N_XI984/QB_XI984/MM4_d N_XI984/Q_XI984/MM4_g N_VDD_XI984/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1035/MM8 N_XI1035/NET08_XI1035/MM8_d N_RWL<15>_XI1035/MM8_g
+ N_RBL<1>_XI1035/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1035/MM7 N_XI1035/NET08_XI1035/MM7_d N_XI1035/QB_XI1035/MM7_g
+ N_GND_XI1035/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1035/MM10 N_WBL<1>_XI1035/MM10_d N_WWLB<15>_XI1035/MM10_g
+ N_XI1035/Q_XI1035/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1035/MM11 N_WBLB<1>_XI1035/MM11_d N_WWLB<15>_XI1035/MM11_g
+ N_XI1035/QB_XI1035/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1035/MM1 N_XI1035/Q_XI1035/MM1_d N_XI1035/QB_XI1035/MM1_g N_GND_XI1035/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1035/MM0 N_XI1035/QB_XI1035/MM0_d N_XI1035/Q_XI1035/MM0_g N_GND_XI1035/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1035/MM9 N_XI1035/NET08_XI1035/MM9_d N_RWLB<15>_XI1035/MM9_g
+ N_RBL<1>_XI1035/MM9_s N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1035/MM6 N_XI1035/NET08_XI1035/MM6_d N_XI1035/QB_XI1035/MM6_g
+ N_VDD_XI1035/MM6_s N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1035/MM5 N_XI1035/Q_XI1035/MM5_d N_XI1035/QB_XI1035/MM5_g N_VDD_XI1035/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1035/MM4 N_XI1035/QB_XI1035/MM4_d N_XI1035/Q_XI1035/MM4_g N_VDD_XI1035/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI992/MM8 N_XI992/NET08_XI992/MM8_d N_RWL<13>_XI992/MM8_g N_RBL<12>_XI992/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI992/MM7 N_XI992/NET08_XI992/MM7_d N_XI992/QB_XI992/MM7_g N_GND_XI992/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI992/MM10 N_WBL<12>_XI992/MM10_d N_WWLB<13>_XI992/MM10_g
+ N_XI992/Q_XI992/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI992/MM11 N_WBLB<12>_XI992/MM11_d N_WWLB<13>_XI992/MM11_g
+ N_XI992/QB_XI992/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI992/MM1 N_XI992/Q_XI992/MM1_d N_XI992/QB_XI992/MM1_g N_GND_XI992/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI992/MM0 N_XI992/QB_XI992/MM0_d N_XI992/Q_XI992/MM0_g N_GND_XI992/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI992/MM9 N_XI992/NET08_XI992/MM9_d N_RWLB<13>_XI992/MM9_g
+ N_RBL<12>_XI992/MM9_s N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI992/MM6 N_XI992/NET08_XI992/MM6_d N_XI992/QB_XI992/MM6_g N_VDD_XI992/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI992/MM5 N_XI992/Q_XI992/MM5_d N_XI992/QB_XI992/MM5_g N_VDD_XI992/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI992/MM4 N_XI992/QB_XI992/MM4_d N_XI992/Q_XI992/MM4_g N_VDD_XI992/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI951/MM8 N_XI951/NET08_XI951/MM8_d N_RWL<10>_XI951/MM8_g N_RBL<5>_XI951/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI951/MM7 N_XI951/NET08_XI951/MM7_d N_XI951/QB_XI951/MM7_g N_GND_XI951/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI951/MM10 N_WBL<5>_XI951/MM10_d N_WWLB<10>_XI951/MM10_g N_XI951/Q_XI951/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI951/MM11 N_WBLB<5>_XI951/MM11_d N_WWLB<10>_XI951/MM11_g
+ N_XI951/QB_XI951/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI951/MM1 N_XI951/Q_XI951/MM1_d N_XI951/QB_XI951/MM1_g N_GND_XI951/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI951/MM0 N_XI951/QB_XI951/MM0_d N_XI951/Q_XI951/MM0_g N_GND_XI951/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI951/MM9 N_XI951/NET08_XI951/MM9_d N_RWLB<10>_XI951/MM9_g N_RBL<5>_XI951/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI951/MM6 N_XI951/NET08_XI951/MM6_d N_XI951/QB_XI951/MM6_g N_VDD_XI951/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI951/MM5 N_XI951/Q_XI951/MM5_d N_XI951/QB_XI951/MM5_g N_VDD_XI951/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI951/MM4 N_XI951/QB_XI951/MM4_d N_XI951/Q_XI951/MM4_g N_VDD_XI951/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI950/MM8 N_XI950/NET08_XI950/MM8_d N_RWL<10>_XI950/MM8_g N_RBL<6>_XI950/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI950/MM7 N_XI950/NET08_XI950/MM7_d N_XI950/QB_XI950/MM7_g N_GND_XI950/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI950/MM10 N_WBL<6>_XI950/MM10_d N_WWLB<10>_XI950/MM10_g N_XI950/Q_XI950/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI950/MM11 N_WBLB<6>_XI950/MM11_d N_WWLB<10>_XI950/MM11_g
+ N_XI950/QB_XI950/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI950/MM1 N_XI950/Q_XI950/MM1_d N_XI950/QB_XI950/MM1_g N_GND_XI950/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI950/MM0 N_XI950/QB_XI950/MM0_d N_XI950/Q_XI950/MM0_g N_GND_XI950/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI950/MM9 N_XI950/NET08_XI950/MM9_d N_RWLB<10>_XI950/MM9_g N_RBL<6>_XI950/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI950/MM6 N_XI950/NET08_XI950/MM6_d N_XI950/QB_XI950/MM6_g N_VDD_XI950/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI950/MM5 N_XI950/Q_XI950/MM5_d N_XI950/QB_XI950/MM5_g N_VDD_XI950/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI950/MM4 N_XI950/QB_XI950/MM4_d N_XI950/Q_XI950/MM4_g N_VDD_XI950/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI949/MM8 N_XI949/NET08_XI949/MM8_d N_RWL<10>_XI949/MM8_g N_RBL<7>_XI949/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI949/MM7 N_XI949/NET08_XI949/MM7_d N_XI949/QB_XI949/MM7_g N_GND_XI949/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI949/MM10 N_WBL<7>_XI949/MM10_d N_WWLB<10>_XI949/MM10_g N_XI949/Q_XI949/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI949/MM11 N_WBLB<7>_XI949/MM11_d N_WWLB<10>_XI949/MM11_g
+ N_XI949/QB_XI949/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI949/MM1 N_XI949/Q_XI949/MM1_d N_XI949/QB_XI949/MM1_g N_GND_XI949/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI949/MM0 N_XI949/QB_XI949/MM0_d N_XI949/Q_XI949/MM0_g N_GND_XI949/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI949/MM9 N_XI949/NET08_XI949/MM9_d N_RWLB<10>_XI949/MM9_g N_RBL<7>_XI949/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI949/MM6 N_XI949/NET08_XI949/MM6_d N_XI949/QB_XI949/MM6_g N_VDD_XI949/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI949/MM5 N_XI949/Q_XI949/MM5_d N_XI949/QB_XI949/MM5_g N_VDD_XI949/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI949/MM4 N_XI949/QB_XI949/MM4_d N_XI949/Q_XI949/MM4_g N_VDD_XI949/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI948/MM8 N_XI948/NET08_XI948/MM8_d N_RWL<10>_XI948/MM8_g N_RBL<8>_XI948/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI948/MM7 N_XI948/NET08_XI948/MM7_d N_XI948/QB_XI948/MM7_g N_GND_XI948/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI948/MM10 N_WBL<8>_XI948/MM10_d N_WWLB<10>_XI948/MM10_g N_XI948/Q_XI948/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI948/MM11 N_WBLB<8>_XI948/MM11_d N_WWLB<10>_XI948/MM11_g
+ N_XI948/QB_XI948/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI948/MM1 N_XI948/Q_XI948/MM1_d N_XI948/QB_XI948/MM1_g N_GND_XI948/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI948/MM0 N_XI948/QB_XI948/MM0_d N_XI948/Q_XI948/MM0_g N_GND_XI948/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI948/MM9 N_XI948/NET08_XI948/MM9_d N_RWLB<10>_XI948/MM9_g N_RBL<8>_XI948/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI948/MM6 N_XI948/NET08_XI948/MM6_d N_XI948/QB_XI948/MM6_g N_VDD_XI948/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI948/MM5 N_XI948/Q_XI948/MM5_d N_XI948/QB_XI948/MM5_g N_VDD_XI948/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI948/MM4 N_XI948/QB_XI948/MM4_d N_XI948/Q_XI948/MM4_g N_VDD_XI948/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI975/MM8 N_XI975/NET08_XI975/MM8_d N_RWL<12>_XI975/MM8_g N_RBL<13>_XI975/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI975/MM7 N_XI975/NET08_XI975/MM7_d N_XI975/QB_XI975/MM7_g N_GND_XI975/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI975/MM10 N_WBL<13>_XI975/MM10_d N_WWLB<12>_XI975/MM10_g
+ N_XI975/Q_XI975/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI975/MM11 N_WBLB<13>_XI975/MM11_d N_WWLB<12>_XI975/MM11_g
+ N_XI975/QB_XI975/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI975/MM1 N_XI975/Q_XI975/MM1_d N_XI975/QB_XI975/MM1_g N_GND_XI975/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI975/MM0 N_XI975/QB_XI975/MM0_d N_XI975/Q_XI975/MM0_g N_GND_XI975/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI975/MM9 N_XI975/NET08_XI975/MM9_d N_RWLB<12>_XI975/MM9_g
+ N_RBL<13>_XI975/MM9_s N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI975/MM6 N_XI975/NET08_XI975/MM6_d N_XI975/QB_XI975/MM6_g N_VDD_XI975/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI975/MM5 N_XI975/Q_XI975/MM5_d N_XI975/QB_XI975/MM5_g N_VDD_XI975/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI975/MM4 N_XI975/QB_XI975/MM4_d N_XI975/Q_XI975/MM4_g N_VDD_XI975/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI974/MM8 N_XI974/NET08_XI974/MM8_d N_RWL<12>_XI974/MM8_g N_RBL<14>_XI974/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI974/MM7 N_XI974/NET08_XI974/MM7_d N_XI974/QB_XI974/MM7_g N_GND_XI974/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI974/MM10 N_WBL<14>_XI974/MM10_d N_WWLB<12>_XI974/MM10_g
+ N_XI974/Q_XI974/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI974/MM11 N_WBLB<14>_XI974/MM11_d N_WWLB<12>_XI974/MM11_g
+ N_XI974/QB_XI974/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI974/MM1 N_XI974/Q_XI974/MM1_d N_XI974/QB_XI974/MM1_g N_GND_XI974/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI974/MM0 N_XI974/QB_XI974/MM0_d N_XI974/Q_XI974/MM0_g N_GND_XI974/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI974/MM9 N_XI974/NET08_XI974/MM9_d N_RWLB<12>_XI974/MM9_g
+ N_RBL<14>_XI974/MM9_s N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI974/MM6 N_XI974/NET08_XI974/MM6_d N_XI974/QB_XI974/MM6_g N_VDD_XI974/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI974/MM5 N_XI974/Q_XI974/MM5_d N_XI974/QB_XI974/MM5_g N_VDD_XI974/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI974/MM4 N_XI974/QB_XI974/MM4_d N_XI974/Q_XI974/MM4_g N_VDD_XI974/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI973/MM8 N_XI973/NET08_XI973/MM8_d N_RWL<11>_XI973/MM8_g N_RBL<15>_XI973/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI973/MM7 N_XI973/NET08_XI973/MM7_d N_XI973/QB_XI973/MM7_g N_GND_XI973/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI973/MM10 N_WBL<15>_XI973/MM10_d N_WWLB<11>_XI973/MM10_g
+ N_XI973/Q_XI973/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI973/MM11 N_WBLB<15>_XI973/MM11_d N_WWLB<11>_XI973/MM11_g
+ N_XI973/QB_XI973/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI973/MM1 N_XI973/Q_XI973/MM1_d N_XI973/QB_XI973/MM1_g N_GND_XI973/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI973/MM0 N_XI973/QB_XI973/MM0_d N_XI973/Q_XI973/MM0_g N_GND_XI973/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI973/MM9 N_XI973/NET08_XI973/MM9_d N_RWLB<11>_XI973/MM9_g
+ N_RBL<15>_XI973/MM9_s N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI973/MM6 N_XI973/NET08_XI973/MM6_d N_XI973/QB_XI973/MM6_g N_VDD_XI973/MM6_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI973/MM5 N_XI973/Q_XI973/MM5_d N_XI973/QB_XI973/MM5_g N_VDD_XI973/MM5_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI973/MM4 N_XI973/QB_XI973/MM4_d N_XI973/Q_XI973/MM4_g N_VDD_XI973/MM4_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI972/MM8 N_XI972/NET08_XI972/MM8_d N_RWL<11>_XI972/MM8_g N_RBL<0>_XI972/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI972/MM7 N_XI972/NET08_XI972/MM7_d N_XI972/QB_XI972/MM7_g N_GND_XI972/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI972/MM10 N_WBL<0>_XI972/MM10_d N_WWLB<11>_XI972/MM10_g N_XI972/Q_XI972/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI972/MM11 N_WBLB<0>_XI972/MM11_d N_WWLB<11>_XI972/MM11_g
+ N_XI972/QB_XI972/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI972/MM1 N_XI972/Q_XI972/MM1_d N_XI972/QB_XI972/MM1_g N_GND_XI972/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI972/MM0 N_XI972/QB_XI972/MM0_d N_XI972/Q_XI972/MM0_g N_GND_XI972/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI972/MM9 N_XI972/NET08_XI972/MM9_d N_RWLB<11>_XI972/MM9_g N_RBL<0>_XI972/MM9_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI972/MM6 N_XI972/NET08_XI972/MM6_d N_XI972/QB_XI972/MM6_g N_VDD_XI972/MM6_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI972/MM5 N_XI972/Q_XI972/MM5_d N_XI972/QB_XI972/MM5_g N_VDD_XI972/MM5_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI972/MM4 N_XI972/QB_XI972/MM4_d N_XI972/Q_XI972/MM4_g N_VDD_XI972/MM4_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI971/MM8 N_XI971/NET08_XI971/MM8_d N_RWL<11>_XI971/MM8_g N_RBL<1>_XI971/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI971/MM7 N_XI971/NET08_XI971/MM7_d N_XI971/QB_XI971/MM7_g N_GND_XI971/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI971/MM10 N_WBL<1>_XI971/MM10_d N_WWLB<11>_XI971/MM10_g N_XI971/Q_XI971/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI971/MM11 N_WBLB<1>_XI971/MM11_d N_WWLB<11>_XI971/MM11_g
+ N_XI971/QB_XI971/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI971/MM1 N_XI971/Q_XI971/MM1_d N_XI971/QB_XI971/MM1_g N_GND_XI971/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI971/MM0 N_XI971/QB_XI971/MM0_d N_XI971/Q_XI971/MM0_g N_GND_XI971/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI971/MM9 N_XI971/NET08_XI971/MM9_d N_RWLB<11>_XI971/MM9_g N_RBL<1>_XI971/MM9_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI971/MM6 N_XI971/NET08_XI971/MM6_d N_XI971/QB_XI971/MM6_g N_VDD_XI971/MM6_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI971/MM5 N_XI971/Q_XI971/MM5_d N_XI971/QB_XI971/MM5_g N_VDD_XI971/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI971/MM4 N_XI971/QB_XI971/MM4_d N_XI971/Q_XI971/MM4_g N_VDD_XI971/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI970/MM8 N_XI970/NET08_XI970/MM8_d N_RWL<11>_XI970/MM8_g N_RBL<2>_XI970/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI970/MM7 N_XI970/NET08_XI970/MM7_d N_XI970/QB_XI970/MM7_g N_GND_XI970/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI970/MM10 N_WBL<2>_XI970/MM10_d N_WWLB<11>_XI970/MM10_g N_XI970/Q_XI970/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI970/MM11 N_WBLB<2>_XI970/MM11_d N_WWLB<11>_XI970/MM11_g
+ N_XI970/QB_XI970/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI970/MM1 N_XI970/Q_XI970/MM1_d N_XI970/QB_XI970/MM1_g N_GND_XI970/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI970/MM0 N_XI970/QB_XI970/MM0_d N_XI970/Q_XI970/MM0_g N_GND_XI970/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI970/MM9 N_XI970/NET08_XI970/MM9_d N_RWLB<11>_XI970/MM9_g N_RBL<2>_XI970/MM9_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI970/MM6 N_XI970/NET08_XI970/MM6_d N_XI970/QB_XI970/MM6_g N_VDD_XI970/MM6_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI970/MM5 N_XI970/Q_XI970/MM5_d N_XI970/QB_XI970/MM5_g N_VDD_XI970/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI970/MM4 N_XI970/QB_XI970/MM4_d N_XI970/Q_XI970/MM4_g N_VDD_XI970/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI990/MM8 N_XI990/NET08_XI990/MM8_d N_RWL<13>_XI990/MM8_g N_RBL<14>_XI990/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI990/MM7 N_XI990/NET08_XI990/MM7_d N_XI990/QB_XI990/MM7_g N_GND_XI990/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI990/MM10 N_WBL<14>_XI990/MM10_d N_WWLB<13>_XI990/MM10_g
+ N_XI990/Q_XI990/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI990/MM11 N_WBLB<14>_XI990/MM11_d N_WWLB<13>_XI990/MM11_g
+ N_XI990/QB_XI990/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI990/MM1 N_XI990/Q_XI990/MM1_d N_XI990/QB_XI990/MM1_g N_GND_XI990/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI990/MM0 N_XI990/QB_XI990/MM0_d N_XI990/Q_XI990/MM0_g N_GND_XI990/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI990/MM9 N_XI990/NET08_XI990/MM9_d N_RWLB<13>_XI990/MM9_g
+ N_RBL<14>_XI990/MM9_s N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI990/MM6 N_XI990/NET08_XI990/MM6_d N_XI990/QB_XI990/MM6_g N_VDD_XI990/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI990/MM5 N_XI990/Q_XI990/MM5_d N_XI990/QB_XI990/MM5_g N_VDD_XI990/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI990/MM4 N_XI990/QB_XI990/MM4_d N_XI990/Q_XI990/MM4_g N_VDD_XI990/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI989/MM8 N_XI989/NET08_XI989/MM8_d N_RWL<12>_XI989/MM8_g N_RBL<15>_XI989/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI989/MM7 N_XI989/NET08_XI989/MM7_d N_XI989/QB_XI989/MM7_g N_GND_XI989/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI989/MM10 N_WBL<15>_XI989/MM10_d N_WWLB<12>_XI989/MM10_g
+ N_XI989/Q_XI989/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI989/MM11 N_WBLB<15>_XI989/MM11_d N_WWLB<12>_XI989/MM11_g
+ N_XI989/QB_XI989/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI989/MM1 N_XI989/Q_XI989/MM1_d N_XI989/QB_XI989/MM1_g N_GND_XI989/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI989/MM0 N_XI989/QB_XI989/MM0_d N_XI989/Q_XI989/MM0_g N_GND_XI989/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI989/MM9 N_XI989/NET08_XI989/MM9_d N_RWLB<12>_XI989/MM9_g
+ N_RBL<15>_XI989/MM9_s N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI989/MM6 N_XI989/NET08_XI989/MM6_d N_XI989/QB_XI989/MM6_g N_VDD_XI989/MM6_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI989/MM5 N_XI989/Q_XI989/MM5_d N_XI989/QB_XI989/MM5_g N_VDD_XI989/MM5_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI989/MM4 N_XI989/QB_XI989/MM4_d N_XI989/Q_XI989/MM4_g N_VDD_XI989/MM4_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI988/MM8 N_XI988/NET08_XI988/MM8_d N_RWL<12>_XI988/MM8_g N_RBL<0>_XI988/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI988/MM7 N_XI988/NET08_XI988/MM7_d N_XI988/QB_XI988/MM7_g N_GND_XI988/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI988/MM10 N_WBL<0>_XI988/MM10_d N_WWLB<12>_XI988/MM10_g N_XI988/Q_XI988/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI988/MM11 N_WBLB<0>_XI988/MM11_d N_WWLB<12>_XI988/MM11_g
+ N_XI988/QB_XI988/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI988/MM1 N_XI988/Q_XI988/MM1_d N_XI988/QB_XI988/MM1_g N_GND_XI988/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI988/MM0 N_XI988/QB_XI988/MM0_d N_XI988/Q_XI988/MM0_g N_GND_XI988/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI988/MM9 N_XI988/NET08_XI988/MM9_d N_RWLB<12>_XI988/MM9_g N_RBL<0>_XI988/MM9_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI988/MM6 N_XI988/NET08_XI988/MM6_d N_XI988/QB_XI988/MM6_g N_VDD_XI988/MM6_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI988/MM5 N_XI988/Q_XI988/MM5_d N_XI988/QB_XI988/MM5_g N_VDD_XI988/MM5_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI988/MM4 N_XI988/QB_XI988/MM4_d N_XI988/Q_XI988/MM4_g N_VDD_XI988/MM4_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI991/MM8 N_XI991/NET08_XI991/MM8_d N_RWL<13>_XI991/MM8_g N_RBL<13>_XI991/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI991/MM7 N_XI991/NET08_XI991/MM7_d N_XI991/QB_XI991/MM7_g N_GND_XI991/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI991/MM10 N_WBL<13>_XI991/MM10_d N_WWLB<13>_XI991/MM10_g
+ N_XI991/Q_XI991/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI991/MM11 N_WBLB<13>_XI991/MM11_d N_WWLB<13>_XI991/MM11_g
+ N_XI991/QB_XI991/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI991/MM1 N_XI991/Q_XI991/MM1_d N_XI991/QB_XI991/MM1_g N_GND_XI991/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI991/MM0 N_XI991/QB_XI991/MM0_d N_XI991/Q_XI991/MM0_g N_GND_XI991/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI991/MM9 N_XI991/NET08_XI991/MM9_d N_RWLB<13>_XI991/MM9_g
+ N_RBL<13>_XI991/MM9_s N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI991/MM6 N_XI991/NET08_XI991/MM6_d N_XI991/QB_XI991/MM6_g N_VDD_XI991/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI991/MM5 N_XI991/Q_XI991/MM5_d N_XI991/QB_XI991/MM5_g N_VDD_XI991/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI991/MM4 N_XI991/QB_XI991/MM4_d N_XI991/Q_XI991/MM4_g N_VDD_XI991/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI981/MM8 N_XI981/NET08_XI981/MM8_d N_RWL<12>_XI981/MM8_g N_RBL<7>_XI981/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI981/MM7 N_XI981/NET08_XI981/MM7_d N_XI981/QB_XI981/MM7_g N_GND_XI981/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI981/MM10 N_WBL<7>_XI981/MM10_d N_WWLB<12>_XI981/MM10_g N_XI981/Q_XI981/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI981/MM11 N_WBLB<7>_XI981/MM11_d N_WWLB<12>_XI981/MM11_g
+ N_XI981/QB_XI981/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI981/MM1 N_XI981/Q_XI981/MM1_d N_XI981/QB_XI981/MM1_g N_GND_XI981/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI981/MM0 N_XI981/QB_XI981/MM0_d N_XI981/Q_XI981/MM0_g N_GND_XI981/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI981/MM9 N_XI981/NET08_XI981/MM9_d N_RWLB<12>_XI981/MM9_g N_RBL<7>_XI981/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI981/MM6 N_XI981/NET08_XI981/MM6_d N_XI981/QB_XI981/MM6_g N_VDD_XI981/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI981/MM5 N_XI981/Q_XI981/MM5_d N_XI981/QB_XI981/MM5_g N_VDD_XI981/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI981/MM4 N_XI981/QB_XI981/MM4_d N_XI981/Q_XI981/MM4_g N_VDD_XI981/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI980/MM8 N_XI980/NET08_XI980/MM8_d N_RWL<12>_XI980/MM8_g N_RBL<8>_XI980/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI980/MM7 N_XI980/NET08_XI980/MM7_d N_XI980/QB_XI980/MM7_g N_GND_XI980/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI980/MM10 N_WBL<8>_XI980/MM10_d N_WWLB<12>_XI980/MM10_g N_XI980/Q_XI980/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI980/MM11 N_WBLB<8>_XI980/MM11_d N_WWLB<12>_XI980/MM11_g
+ N_XI980/QB_XI980/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI980/MM1 N_XI980/Q_XI980/MM1_d N_XI980/QB_XI980/MM1_g N_GND_XI980/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI980/MM0 N_XI980/QB_XI980/MM0_d N_XI980/Q_XI980/MM0_g N_GND_XI980/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI980/MM9 N_XI980/NET08_XI980/MM9_d N_RWLB<12>_XI980/MM9_g N_RBL<8>_XI980/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI980/MM6 N_XI980/NET08_XI980/MM6_d N_XI980/QB_XI980/MM6_g N_VDD_XI980/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI980/MM5 N_XI980/Q_XI980/MM5_d N_XI980/QB_XI980/MM5_g N_VDD_XI980/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI980/MM4 N_XI980/QB_XI980/MM4_d N_XI980/Q_XI980/MM4_g N_VDD_XI980/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1034/MM8 N_XI1034/NET08_XI1034/MM8_d N_RWL<15>_XI1034/MM8_g
+ N_RBL<2>_XI1034/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1034/MM7 N_XI1034/NET08_XI1034/MM7_d N_XI1034/QB_XI1034/MM7_g
+ N_GND_XI1034/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1034/MM10 N_WBL<2>_XI1034/MM10_d N_WWLB<15>_XI1034/MM10_g
+ N_XI1034/Q_XI1034/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1034/MM11 N_WBLB<2>_XI1034/MM11_d N_WWLB<15>_XI1034/MM11_g
+ N_XI1034/QB_XI1034/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1034/MM1 N_XI1034/Q_XI1034/MM1_d N_XI1034/QB_XI1034/MM1_g N_GND_XI1034/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1034/MM0 N_XI1034/QB_XI1034/MM0_d N_XI1034/Q_XI1034/MM0_g N_GND_XI1034/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1034/MM9 N_XI1034/NET08_XI1034/MM9_d N_RWLB<15>_XI1034/MM9_g
+ N_RBL<2>_XI1034/MM9_s N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1034/MM6 N_XI1034/NET08_XI1034/MM6_d N_XI1034/QB_XI1034/MM6_g
+ N_VDD_XI1034/MM6_s N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1034/MM5 N_XI1034/Q_XI1034/MM5_d N_XI1034/QB_XI1034/MM5_g N_VDD_XI1034/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1034/MM4 N_XI1034/QB_XI1034/MM4_d N_XI1034/Q_XI1034/MM4_g N_VDD_XI1034/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI993/MM8 N_XI993/NET08_XI993/MM8_d N_RWL<13>_XI993/MM8_g N_RBL<11>_XI993/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI993/MM7 N_XI993/NET08_XI993/MM7_d N_XI993/QB_XI993/MM7_g N_GND_XI993/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI993/MM10 N_WBL<11>_XI993/MM10_d N_WWLB<13>_XI993/MM10_g
+ N_XI993/Q_XI993/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI993/MM11 N_WBLB<11>_XI993/MM11_d N_WWLB<13>_XI993/MM11_g
+ N_XI993/QB_XI993/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI993/MM1 N_XI993/Q_XI993/MM1_d N_XI993/QB_XI993/MM1_g N_GND_XI993/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI993/MM0 N_XI993/QB_XI993/MM0_d N_XI993/Q_XI993/MM0_g N_GND_XI993/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI993/MM9 N_XI993/NET08_XI993/MM9_d N_RWLB<13>_XI993/MM9_g
+ N_RBL<11>_XI993/MM9_s N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI993/MM6 N_XI993/NET08_XI993/MM6_d N_XI993/QB_XI993/MM6_g N_VDD_XI993/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI993/MM5 N_XI993/Q_XI993/MM5_d N_XI993/QB_XI993/MM5_g N_VDD_XI993/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI993/MM4 N_XI993/QB_XI993/MM4_d N_XI993/Q_XI993/MM4_g N_VDD_XI993/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI947/MM8 N_XI947/NET08_XI947/MM8_d N_RWL<10>_XI947/MM8_g N_RBL<9>_XI947/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI947/MM7 N_XI947/NET08_XI947/MM7_d N_XI947/QB_XI947/MM7_g N_GND_XI947/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI947/MM10 N_WBL<9>_XI947/MM10_d N_WWLB<10>_XI947/MM10_g N_XI947/Q_XI947/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI947/MM11 N_WBLB<9>_XI947/MM11_d N_WWLB<10>_XI947/MM11_g
+ N_XI947/QB_XI947/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI947/MM1 N_XI947/Q_XI947/MM1_d N_XI947/QB_XI947/MM1_g N_GND_XI947/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI947/MM0 N_XI947/QB_XI947/MM0_d N_XI947/Q_XI947/MM0_g N_GND_XI947/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI947/MM9 N_XI947/NET08_XI947/MM9_d N_RWLB<10>_XI947/MM9_g N_RBL<9>_XI947/MM9_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI947/MM6 N_XI947/NET08_XI947/MM6_d N_XI947/QB_XI947/MM6_g N_VDD_XI947/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI947/MM5 N_XI947/Q_XI947/MM5_d N_XI947/QB_XI947/MM5_g N_VDD_XI947/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI947/MM4 N_XI947/QB_XI947/MM4_d N_XI947/Q_XI947/MM4_g N_VDD_XI947/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI946/MM8 N_XI946/NET08_XI946/MM8_d N_RWL<10>_XI946/MM8_g N_RBL<10>_XI946/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI946/MM7 N_XI946/NET08_XI946/MM7_d N_XI946/QB_XI946/MM7_g N_GND_XI946/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI946/MM10 N_WBL<10>_XI946/MM10_d N_WWLB<10>_XI946/MM10_g
+ N_XI946/Q_XI946/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI946/MM11 N_WBLB<10>_XI946/MM11_d N_WWLB<10>_XI946/MM11_g
+ N_XI946/QB_XI946/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI946/MM1 N_XI946/Q_XI946/MM1_d N_XI946/QB_XI946/MM1_g N_GND_XI946/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI946/MM0 N_XI946/QB_XI946/MM0_d N_XI946/Q_XI946/MM0_g N_GND_XI946/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI946/MM9 N_XI946/NET08_XI946/MM9_d N_RWLB<10>_XI946/MM9_g
+ N_RBL<10>_XI946/MM9_s N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI946/MM6 N_XI946/NET08_XI946/MM6_d N_XI946/QB_XI946/MM6_g N_VDD_XI946/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI946/MM5 N_XI946/Q_XI946/MM5_d N_XI946/QB_XI946/MM5_g N_VDD_XI946/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI946/MM4 N_XI946/QB_XI946/MM4_d N_XI946/Q_XI946/MM4_g N_VDD_XI946/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI945/MM8 N_XI945/NET08_XI945/MM8_d N_RWL<10>_XI945/MM8_g N_RBL<11>_XI945/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI945/MM7 N_XI945/NET08_XI945/MM7_d N_XI945/QB_XI945/MM7_g N_GND_XI945/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI945/MM10 N_WBL<11>_XI945/MM10_d N_WWLB<10>_XI945/MM10_g
+ N_XI945/Q_XI945/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI945/MM11 N_WBLB<11>_XI945/MM11_d N_WWLB<10>_XI945/MM11_g
+ N_XI945/QB_XI945/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI945/MM1 N_XI945/Q_XI945/MM1_d N_XI945/QB_XI945/MM1_g N_GND_XI945/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI945/MM0 N_XI945/QB_XI945/MM0_d N_XI945/Q_XI945/MM0_g N_GND_XI945/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI945/MM9 N_XI945/NET08_XI945/MM9_d N_RWLB<10>_XI945/MM9_g
+ N_RBL<11>_XI945/MM9_s N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI945/MM6 N_XI945/NET08_XI945/MM6_d N_XI945/QB_XI945/MM6_g N_VDD_XI945/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI945/MM5 N_XI945/Q_XI945/MM5_d N_XI945/QB_XI945/MM5_g N_VDD_XI945/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI945/MM4 N_XI945/QB_XI945/MM4_d N_XI945/Q_XI945/MM4_g N_VDD_XI945/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI944/MM8 N_XI944/NET08_XI944/MM8_d N_RWL<10>_XI944/MM8_g N_RBL<12>_XI944/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI944/MM7 N_XI944/NET08_XI944/MM7_d N_XI944/QB_XI944/MM7_g N_GND_XI944/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI944/MM10 N_WBL<12>_XI944/MM10_d N_WWLB<10>_XI944/MM10_g
+ N_XI944/Q_XI944/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI944/MM11 N_WBLB<12>_XI944/MM11_d N_WWLB<10>_XI944/MM11_g
+ N_XI944/QB_XI944/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI944/MM1 N_XI944/Q_XI944/MM1_d N_XI944/QB_XI944/MM1_g N_GND_XI944/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI944/MM0 N_XI944/QB_XI944/MM0_d N_XI944/Q_XI944/MM0_g N_GND_XI944/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI944/MM9 N_XI944/NET08_XI944/MM9_d N_RWLB<10>_XI944/MM9_g
+ N_RBL<12>_XI944/MM9_s N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI944/MM6 N_XI944/NET08_XI944/MM6_d N_XI944/QB_XI944/MM6_g N_VDD_XI944/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI944/MM5 N_XI944/Q_XI944/MM5_d N_XI944/QB_XI944/MM5_g N_VDD_XI944/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI944/MM4 N_XI944/QB_XI944/MM4_d N_XI944/Q_XI944/MM4_g N_VDD_XI944/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI969/MM8 N_XI969/NET08_XI969/MM8_d N_RWL<11>_XI969/MM8_g N_RBL<3>_XI969/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI969/MM7 N_XI969/NET08_XI969/MM7_d N_XI969/QB_XI969/MM7_g N_GND_XI969/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI969/MM10 N_WBL<3>_XI969/MM10_d N_WWLB<11>_XI969/MM10_g N_XI969/Q_XI969/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI969/MM11 N_WBLB<3>_XI969/MM11_d N_WWLB<11>_XI969/MM11_g
+ N_XI969/QB_XI969/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI969/MM1 N_XI969/Q_XI969/MM1_d N_XI969/QB_XI969/MM1_g N_GND_XI969/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI969/MM0 N_XI969/QB_XI969/MM0_d N_XI969/Q_XI969/MM0_g N_GND_XI969/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI969/MM9 N_XI969/NET08_XI969/MM9_d N_RWLB<11>_XI969/MM9_g N_RBL<3>_XI969/MM9_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI969/MM6 N_XI969/NET08_XI969/MM6_d N_XI969/QB_XI969/MM6_g N_VDD_XI969/MM6_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI969/MM5 N_XI969/Q_XI969/MM5_d N_XI969/QB_XI969/MM5_g N_VDD_XI969/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI969/MM4 N_XI969/QB_XI969/MM4_d N_XI969/Q_XI969/MM4_g N_VDD_XI969/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI968/MM8 N_XI968/NET08_XI968/MM8_d N_RWL<11>_XI968/MM8_g N_RBL<4>_XI968/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI968/MM7 N_XI968/NET08_XI968/MM7_d N_XI968/QB_XI968/MM7_g N_GND_XI968/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI968/MM10 N_WBL<4>_XI968/MM10_d N_WWLB<11>_XI968/MM10_g N_XI968/Q_XI968/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI968/MM11 N_WBLB<4>_XI968/MM11_d N_WWLB<11>_XI968/MM11_g
+ N_XI968/QB_XI968/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI968/MM1 N_XI968/Q_XI968/MM1_d N_XI968/QB_XI968/MM1_g N_GND_XI968/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI968/MM0 N_XI968/QB_XI968/MM0_d N_XI968/Q_XI968/MM0_g N_GND_XI968/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI968/MM9 N_XI968/NET08_XI968/MM9_d N_RWLB<11>_XI968/MM9_g N_RBL<4>_XI968/MM9_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI968/MM6 N_XI968/NET08_XI968/MM6_d N_XI968/QB_XI968/MM6_g N_VDD_XI968/MM6_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI968/MM5 N_XI968/Q_XI968/MM5_d N_XI968/QB_XI968/MM5_g N_VDD_XI968/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI968/MM4 N_XI968/QB_XI968/MM4_d N_XI968/Q_XI968/MM4_g N_VDD_XI968/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI967/MM8 N_XI967/NET08_XI967/MM8_d N_RWL<11>_XI967/MM8_g N_RBL<5>_XI967/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI967/MM7 N_XI967/NET08_XI967/MM7_d N_XI967/QB_XI967/MM7_g N_GND_XI967/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI967/MM10 N_WBL<5>_XI967/MM10_d N_WWLB<11>_XI967/MM10_g N_XI967/Q_XI967/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI967/MM11 N_WBLB<5>_XI967/MM11_d N_WWLB<11>_XI967/MM11_g
+ N_XI967/QB_XI967/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI967/MM1 N_XI967/Q_XI967/MM1_d N_XI967/QB_XI967/MM1_g N_GND_XI967/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI967/MM0 N_XI967/QB_XI967/MM0_d N_XI967/Q_XI967/MM0_g N_GND_XI967/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI967/MM9 N_XI967/NET08_XI967/MM9_d N_RWLB<11>_XI967/MM9_g N_RBL<5>_XI967/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI967/MM6 N_XI967/NET08_XI967/MM6_d N_XI967/QB_XI967/MM6_g N_VDD_XI967/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI967/MM5 N_XI967/Q_XI967/MM5_d N_XI967/QB_XI967/MM5_g N_VDD_XI967/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI967/MM4 N_XI967/QB_XI967/MM4_d N_XI967/Q_XI967/MM4_g N_VDD_XI967/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI966/MM8 N_XI966/NET08_XI966/MM8_d N_RWL<11>_XI966/MM8_g N_RBL<6>_XI966/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI966/MM7 N_XI966/NET08_XI966/MM7_d N_XI966/QB_XI966/MM7_g N_GND_XI966/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI966/MM10 N_WBL<6>_XI966/MM10_d N_WWLB<11>_XI966/MM10_g N_XI966/Q_XI966/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI966/MM11 N_WBLB<6>_XI966/MM11_d N_WWLB<11>_XI966/MM11_g
+ N_XI966/QB_XI966/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI966/MM1 N_XI966/Q_XI966/MM1_d N_XI966/QB_XI966/MM1_g N_GND_XI966/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI966/MM0 N_XI966/QB_XI966/MM0_d N_XI966/Q_XI966/MM0_g N_GND_XI966/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI966/MM9 N_XI966/NET08_XI966/MM9_d N_RWLB<11>_XI966/MM9_g N_RBL<6>_XI966/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI966/MM6 N_XI966/NET08_XI966/MM6_d N_XI966/QB_XI966/MM6_g N_VDD_XI966/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI966/MM5 N_XI966/Q_XI966/MM5_d N_XI966/QB_XI966/MM5_g N_VDD_XI966/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI966/MM4 N_XI966/QB_XI966/MM4_d N_XI966/Q_XI966/MM4_g N_VDD_XI966/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI965/MM8 N_XI965/NET08_XI965/MM8_d N_RWL<11>_XI965/MM8_g N_RBL<7>_XI965/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI965/MM7 N_XI965/NET08_XI965/MM7_d N_XI965/QB_XI965/MM7_g N_GND_XI965/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI965/MM10 N_WBL<7>_XI965/MM10_d N_WWLB<11>_XI965/MM10_g N_XI965/Q_XI965/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI965/MM11 N_WBLB<7>_XI965/MM11_d N_WWLB<11>_XI965/MM11_g
+ N_XI965/QB_XI965/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI965/MM1 N_XI965/Q_XI965/MM1_d N_XI965/QB_XI965/MM1_g N_GND_XI965/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI965/MM0 N_XI965/QB_XI965/MM0_d N_XI965/Q_XI965/MM0_g N_GND_XI965/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI965/MM9 N_XI965/NET08_XI965/MM9_d N_RWLB<11>_XI965/MM9_g N_RBL<7>_XI965/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI965/MM6 N_XI965/NET08_XI965/MM6_d N_XI965/QB_XI965/MM6_g N_VDD_XI965/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI965/MM5 N_XI965/Q_XI965/MM5_d N_XI965/QB_XI965/MM5_g N_VDD_XI965/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI965/MM4 N_XI965/QB_XI965/MM4_d N_XI965/Q_XI965/MM4_g N_VDD_XI965/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI964/MM8 N_XI964/NET08_XI964/MM8_d N_RWL<11>_XI964/MM8_g N_RBL<8>_XI964/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI964/MM7 N_XI964/NET08_XI964/MM7_d N_XI964/QB_XI964/MM7_g N_GND_XI964/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI964/MM10 N_WBL<8>_XI964/MM10_d N_WWLB<11>_XI964/MM10_g N_XI964/Q_XI964/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI964/MM11 N_WBLB<8>_XI964/MM11_d N_WWLB<11>_XI964/MM11_g
+ N_XI964/QB_XI964/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI964/MM1 N_XI964/Q_XI964/MM1_d N_XI964/QB_XI964/MM1_g N_GND_XI964/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI964/MM0 N_XI964/QB_XI964/MM0_d N_XI964/Q_XI964/MM0_g N_GND_XI964/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI964/MM9 N_XI964/NET08_XI964/MM9_d N_RWLB<11>_XI964/MM9_g N_RBL<8>_XI964/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI964/MM6 N_XI964/NET08_XI964/MM6_d N_XI964/QB_XI964/MM6_g N_VDD_XI964/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI964/MM5 N_XI964/Q_XI964/MM5_d N_XI964/QB_XI964/MM5_g N_VDD_XI964/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI964/MM4 N_XI964/QB_XI964/MM4_d N_XI964/Q_XI964/MM4_g N_VDD_XI964/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI987/MM8 N_XI987/NET08_XI987/MM8_d N_RWL<12>_XI987/MM8_g N_RBL<1>_XI987/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI987/MM7 N_XI987/NET08_XI987/MM7_d N_XI987/QB_XI987/MM7_g N_GND_XI987/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI987/MM10 N_WBL<1>_XI987/MM10_d N_WWLB<12>_XI987/MM10_g N_XI987/Q_XI987/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI987/MM11 N_WBLB<1>_XI987/MM11_d N_WWLB<12>_XI987/MM11_g
+ N_XI987/QB_XI987/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI987/MM1 N_XI987/Q_XI987/MM1_d N_XI987/QB_XI987/MM1_g N_GND_XI987/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI987/MM0 N_XI987/QB_XI987/MM0_d N_XI987/Q_XI987/MM0_g N_GND_XI987/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI987/MM9 N_XI987/NET08_XI987/MM9_d N_RWLB<12>_XI987/MM9_g N_RBL<1>_XI987/MM9_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI987/MM6 N_XI987/NET08_XI987/MM6_d N_XI987/QB_XI987/MM6_g N_VDD_XI987/MM6_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI987/MM5 N_XI987/Q_XI987/MM5_d N_XI987/QB_XI987/MM5_g N_VDD_XI987/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI987/MM4 N_XI987/QB_XI987/MM4_d N_XI987/Q_XI987/MM4_g N_VDD_XI987/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI986/MM8 N_XI986/NET08_XI986/MM8_d N_RWL<12>_XI986/MM8_g N_RBL<2>_XI986/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI986/MM7 N_XI986/NET08_XI986/MM7_d N_XI986/QB_XI986/MM7_g N_GND_XI986/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI986/MM10 N_WBL<2>_XI986/MM10_d N_WWLB<12>_XI986/MM10_g N_XI986/Q_XI986/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI986/MM11 N_WBLB<2>_XI986/MM11_d N_WWLB<12>_XI986/MM11_g
+ N_XI986/QB_XI986/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI986/MM1 N_XI986/Q_XI986/MM1_d N_XI986/QB_XI986/MM1_g N_GND_XI986/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI986/MM0 N_XI986/QB_XI986/MM0_d N_XI986/Q_XI986/MM0_g N_GND_XI986/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI986/MM9 N_XI986/NET08_XI986/MM9_d N_RWLB<12>_XI986/MM9_g N_RBL<2>_XI986/MM9_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI986/MM6 N_XI986/NET08_XI986/MM6_d N_XI986/QB_XI986/MM6_g N_VDD_XI986/MM6_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI986/MM5 N_XI986/Q_XI986/MM5_d N_XI986/QB_XI986/MM5_g N_VDD_XI986/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI986/MM4 N_XI986/QB_XI986/MM4_d N_XI986/Q_XI986/MM4_g N_VDD_XI986/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI985/MM8 N_XI985/NET08_XI985/MM8_d N_RWL<12>_XI985/MM8_g N_RBL<3>_XI985/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI985/MM7 N_XI985/NET08_XI985/MM7_d N_XI985/QB_XI985/MM7_g N_GND_XI985/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI985/MM10 N_WBL<3>_XI985/MM10_d N_WWLB<12>_XI985/MM10_g N_XI985/Q_XI985/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI985/MM11 N_WBLB<3>_XI985/MM11_d N_WWLB<12>_XI985/MM11_g
+ N_XI985/QB_XI985/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI985/MM1 N_XI985/Q_XI985/MM1_d N_XI985/QB_XI985/MM1_g N_GND_XI985/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI985/MM0 N_XI985/QB_XI985/MM0_d N_XI985/Q_XI985/MM0_g N_GND_XI985/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI985/MM9 N_XI985/NET08_XI985/MM9_d N_RWLB<12>_XI985/MM9_g N_RBL<3>_XI985/MM9_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI985/MM6 N_XI985/NET08_XI985/MM6_d N_XI985/QB_XI985/MM6_g N_VDD_XI985/MM6_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI985/MM5 N_XI985/Q_XI985/MM5_d N_XI985/QB_XI985/MM5_g N_VDD_XI985/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI985/MM4 N_XI985/QB_XI985/MM4_d N_XI985/Q_XI985/MM4_g N_VDD_XI985/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI978/MM8 N_XI978/NET08_XI978/MM8_d N_RWL<12>_XI978/MM8_g N_RBL<10>_XI978/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI978/MM7 N_XI978/NET08_XI978/MM7_d N_XI978/QB_XI978/MM7_g N_GND_XI978/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI978/MM10 N_WBL<10>_XI978/MM10_d N_WWLB<12>_XI978/MM10_g
+ N_XI978/Q_XI978/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI978/MM11 N_WBLB<10>_XI978/MM11_d N_WWLB<12>_XI978/MM11_g
+ N_XI978/QB_XI978/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI978/MM1 N_XI978/Q_XI978/MM1_d N_XI978/QB_XI978/MM1_g N_GND_XI978/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI978/MM0 N_XI978/QB_XI978/MM0_d N_XI978/Q_XI978/MM0_g N_GND_XI978/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI978/MM9 N_XI978/NET08_XI978/MM9_d N_RWLB<12>_XI978/MM9_g
+ N_RBL<10>_XI978/MM9_s N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI978/MM6 N_XI978/NET08_XI978/MM6_d N_XI978/QB_XI978/MM6_g N_VDD_XI978/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI978/MM5 N_XI978/Q_XI978/MM5_d N_XI978/QB_XI978/MM5_g N_VDD_XI978/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI978/MM4 N_XI978/QB_XI978/MM4_d N_XI978/Q_XI978/MM4_g N_VDD_XI978/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI977/MM8 N_XI977/NET08_XI977/MM8_d N_RWL<12>_XI977/MM8_g N_RBL<11>_XI977/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI977/MM7 N_XI977/NET08_XI977/MM7_d N_XI977/QB_XI977/MM7_g N_GND_XI977/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI977/MM10 N_WBL<11>_XI977/MM10_d N_WWLB<12>_XI977/MM10_g
+ N_XI977/Q_XI977/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI977/MM11 N_WBLB<11>_XI977/MM11_d N_WWLB<12>_XI977/MM11_g
+ N_XI977/QB_XI977/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI977/MM1 N_XI977/Q_XI977/MM1_d N_XI977/QB_XI977/MM1_g N_GND_XI977/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI977/MM0 N_XI977/QB_XI977/MM0_d N_XI977/Q_XI977/MM0_g N_GND_XI977/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI977/MM9 N_XI977/NET08_XI977/MM9_d N_RWLB<12>_XI977/MM9_g
+ N_RBL<11>_XI977/MM9_s N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI977/MM6 N_XI977/NET08_XI977/MM6_d N_XI977/QB_XI977/MM6_g N_VDD_XI977/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI977/MM5 N_XI977/Q_XI977/MM5_d N_XI977/QB_XI977/MM5_g N_VDD_XI977/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI977/MM4 N_XI977/QB_XI977/MM4_d N_XI977/Q_XI977/MM4_g N_VDD_XI977/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI976/MM8 N_XI976/NET08_XI976/MM8_d N_RWL<12>_XI976/MM8_g N_RBL<12>_XI976/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI976/MM7 N_XI976/NET08_XI976/MM7_d N_XI976/QB_XI976/MM7_g N_GND_XI976/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI976/MM10 N_WBL<12>_XI976/MM10_d N_WWLB<12>_XI976/MM10_g
+ N_XI976/Q_XI976/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI976/MM11 N_WBLB<12>_XI976/MM11_d N_WWLB<12>_XI976/MM11_g
+ N_XI976/QB_XI976/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI976/MM1 N_XI976/Q_XI976/MM1_d N_XI976/QB_XI976/MM1_g N_GND_XI976/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI976/MM0 N_XI976/QB_XI976/MM0_d N_XI976/Q_XI976/MM0_g N_GND_XI976/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI976/MM9 N_XI976/NET08_XI976/MM9_d N_RWLB<12>_XI976/MM9_g
+ N_RBL<12>_XI976/MM9_s N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI976/MM6 N_XI976/NET08_XI976/MM6_d N_XI976/QB_XI976/MM6_g N_VDD_XI976/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI976/MM5 N_XI976/Q_XI976/MM5_d N_XI976/QB_XI976/MM5_g N_VDD_XI976/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI976/MM4 N_XI976/QB_XI976/MM4_d N_XI976/Q_XI976/MM4_g N_VDD_XI976/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1033/MM8 N_XI1033/NET08_XI1033/MM8_d N_RWL<15>_XI1033/MM8_g
+ N_RBL<3>_XI1033/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1033/MM7 N_XI1033/NET08_XI1033/MM7_d N_XI1033/QB_XI1033/MM7_g
+ N_GND_XI1033/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1033/MM10 N_WBL<3>_XI1033/MM10_d N_WWLB<15>_XI1033/MM10_g
+ N_XI1033/Q_XI1033/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1033/MM11 N_WBLB<3>_XI1033/MM11_d N_WWLB<15>_XI1033/MM11_g
+ N_XI1033/QB_XI1033/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1033/MM1 N_XI1033/Q_XI1033/MM1_d N_XI1033/QB_XI1033/MM1_g N_GND_XI1033/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1033/MM0 N_XI1033/QB_XI1033/MM0_d N_XI1033/Q_XI1033/MM0_g N_GND_XI1033/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1033/MM9 N_XI1033/NET08_XI1033/MM9_d N_RWLB<15>_XI1033/MM9_g
+ N_RBL<3>_XI1033/MM9_s N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1033/MM6 N_XI1033/NET08_XI1033/MM6_d N_XI1033/QB_XI1033/MM6_g
+ N_VDD_XI1033/MM6_s N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1033/MM5 N_XI1033/Q_XI1033/MM5_d N_XI1033/QB_XI1033/MM5_g N_VDD_XI1033/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1033/MM4 N_XI1033/QB_XI1033/MM4_d N_XI1033/Q_XI1033/MM4_g N_VDD_XI1033/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI994/MM8 N_XI994/NET08_XI994/MM8_d N_RWL<13>_XI994/MM8_g N_RBL<10>_XI994/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI994/MM7 N_XI994/NET08_XI994/MM7_d N_XI994/QB_XI994/MM7_g N_GND_XI994/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI994/MM10 N_WBL<10>_XI994/MM10_d N_WWLB<13>_XI994/MM10_g
+ N_XI994/Q_XI994/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI994/MM11 N_WBLB<10>_XI994/MM11_d N_WWLB<13>_XI994/MM11_g
+ N_XI994/QB_XI994/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI994/MM1 N_XI994/Q_XI994/MM1_d N_XI994/QB_XI994/MM1_g N_GND_XI994/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI994/MM0 N_XI994/QB_XI994/MM0_d N_XI994/Q_XI994/MM0_g N_GND_XI994/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI994/MM9 N_XI994/NET08_XI994/MM9_d N_RWLB<13>_XI994/MM9_g
+ N_RBL<10>_XI994/MM9_s N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI994/MM6 N_XI994/NET08_XI994/MM6_d N_XI994/QB_XI994/MM6_g N_VDD_XI994/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI994/MM5 N_XI994/Q_XI994/MM5_d N_XI994/QB_XI994/MM5_g N_VDD_XI994/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI994/MM4 N_XI994/QB_XI994/MM4_d N_XI994/Q_XI994/MM4_g N_VDD_XI994/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI943/MM8 N_XI943/NET08_XI943/MM8_d N_RWL<10>_XI943/MM8_g N_RBL<13>_XI943/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI943/MM7 N_XI943/NET08_XI943/MM7_d N_XI943/QB_XI943/MM7_g N_GND_XI943/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI943/MM10 N_WBL<13>_XI943/MM10_d N_WWLB<10>_XI943/MM10_g
+ N_XI943/Q_XI943/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI943/MM11 N_WBLB<13>_XI943/MM11_d N_WWLB<10>_XI943/MM11_g
+ N_XI943/QB_XI943/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI943/MM1 N_XI943/Q_XI943/MM1_d N_XI943/QB_XI943/MM1_g N_GND_XI943/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI943/MM0 N_XI943/QB_XI943/MM0_d N_XI943/Q_XI943/MM0_g N_GND_XI943/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI943/MM9 N_XI943/NET08_XI943/MM9_d N_RWLB<10>_XI943/MM9_g
+ N_RBL<13>_XI943/MM9_s N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI943/MM6 N_XI943/NET08_XI943/MM6_d N_XI943/QB_XI943/MM6_g N_VDD_XI943/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI943/MM5 N_XI943/Q_XI943/MM5_d N_XI943/QB_XI943/MM5_g N_VDD_XI943/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI943/MM4 N_XI943/QB_XI943/MM4_d N_XI943/Q_XI943/MM4_g N_VDD_XI943/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI942/MM8 N_XI942/NET08_XI942/MM8_d N_RWL<10>_XI942/MM8_g N_RBL<14>_XI942/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI942/MM7 N_XI942/NET08_XI942/MM7_d N_XI942/QB_XI942/MM7_g N_GND_XI942/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI942/MM10 N_WBL<14>_XI942/MM10_d N_WWLB<10>_XI942/MM10_g
+ N_XI942/Q_XI942/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI942/MM11 N_WBLB<14>_XI942/MM11_d N_WWLB<10>_XI942/MM11_g
+ N_XI942/QB_XI942/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI942/MM1 N_XI942/Q_XI942/MM1_d N_XI942/QB_XI942/MM1_g N_GND_XI942/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI942/MM0 N_XI942/QB_XI942/MM0_d N_XI942/Q_XI942/MM0_g N_GND_XI942/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI942/MM9 N_XI942/NET08_XI942/MM9_d N_RWLB<10>_XI942/MM9_g
+ N_RBL<14>_XI942/MM9_s N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI942/MM6 N_XI942/NET08_XI942/MM6_d N_XI942/QB_XI942/MM6_g N_VDD_XI942/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI942/MM5 N_XI942/Q_XI942/MM5_d N_XI942/QB_XI942/MM5_g N_VDD_XI942/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI942/MM4 N_XI942/QB_XI942/MM4_d N_XI942/Q_XI942/MM4_g N_VDD_XI942/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI941/MM8 N_XI941/NET08_XI941/MM8_d N_RWL<9>_XI941/MM8_g N_RBL<15>_XI941/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI941/MM7 N_XI941/NET08_XI941/MM7_d N_XI941/QB_XI941/MM7_g N_GND_XI941/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI941/MM10 N_WBL<15>_XI941/MM10_d N_WWLB<9>_XI941/MM10_g N_XI941/Q_XI941/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI941/MM11 N_WBLB<15>_XI941/MM11_d N_WWLB<9>_XI941/MM11_g
+ N_XI941/QB_XI941/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI941/MM1 N_XI941/Q_XI941/MM1_d N_XI941/QB_XI941/MM1_g N_GND_XI941/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI941/MM0 N_XI941/QB_XI941/MM0_d N_XI941/Q_XI941/MM0_g N_GND_XI941/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI941/MM9 N_XI941/NET08_XI941/MM9_d N_RWLB<9>_XI941/MM9_g N_RBL<15>_XI941/MM9_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI941/MM6 N_XI941/NET08_XI941/MM6_d N_XI941/QB_XI941/MM6_g N_VDD_XI941/MM6_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI941/MM5 N_XI941/Q_XI941/MM5_d N_XI941/QB_XI941/MM5_g N_VDD_XI941/MM5_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI941/MM4 N_XI941/QB_XI941/MM4_d N_XI941/Q_XI941/MM4_g N_VDD_XI941/MM4_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI940/MM8 N_XI940/NET08_XI940/MM8_d N_RWL<9>_XI940/MM8_g N_RBL<0>_XI940/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI940/MM7 N_XI940/NET08_XI940/MM7_d N_XI940/QB_XI940/MM7_g N_GND_XI940/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI940/MM10 N_WBL<0>_XI940/MM10_d N_WWLB<9>_XI940/MM10_g N_XI940/Q_XI940/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI940/MM11 N_WBLB<0>_XI940/MM11_d N_WWLB<9>_XI940/MM11_g
+ N_XI940/QB_XI940/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI940/MM1 N_XI940/Q_XI940/MM1_d N_XI940/QB_XI940/MM1_g N_GND_XI940/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI940/MM0 N_XI940/QB_XI940/MM0_d N_XI940/Q_XI940/MM0_g N_GND_XI940/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI940/MM9 N_XI940/NET08_XI940/MM9_d N_RWLB<9>_XI940/MM9_g N_RBL<0>_XI940/MM9_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI940/MM6 N_XI940/NET08_XI940/MM6_d N_XI940/QB_XI940/MM6_g N_VDD_XI940/MM6_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI940/MM5 N_XI940/Q_XI940/MM5_d N_XI940/QB_XI940/MM5_g N_VDD_XI940/MM5_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI940/MM4 N_XI940/QB_XI940/MM4_d N_XI940/Q_XI940/MM4_g N_VDD_XI940/MM4_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI963/MM8 N_XI963/NET08_XI963/MM8_d N_RWL<11>_XI963/MM8_g N_RBL<9>_XI963/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI963/MM7 N_XI963/NET08_XI963/MM7_d N_XI963/QB_XI963/MM7_g N_GND_XI963/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI963/MM10 N_WBL<9>_XI963/MM10_d N_WWLB<11>_XI963/MM10_g N_XI963/Q_XI963/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI963/MM11 N_WBLB<9>_XI963/MM11_d N_WWLB<11>_XI963/MM11_g
+ N_XI963/QB_XI963/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI963/MM1 N_XI963/Q_XI963/MM1_d N_XI963/QB_XI963/MM1_g N_GND_XI963/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI963/MM0 N_XI963/QB_XI963/MM0_d N_XI963/Q_XI963/MM0_g N_GND_XI963/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI963/MM9 N_XI963/NET08_XI963/MM9_d N_RWLB<11>_XI963/MM9_g N_RBL<9>_XI963/MM9_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI963/MM6 N_XI963/NET08_XI963/MM6_d N_XI963/QB_XI963/MM6_g N_VDD_XI963/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI963/MM5 N_XI963/Q_XI963/MM5_d N_XI963/QB_XI963/MM5_g N_VDD_XI963/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI963/MM4 N_XI963/QB_XI963/MM4_d N_XI963/Q_XI963/MM4_g N_VDD_XI963/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI962/MM8 N_XI962/NET08_XI962/MM8_d N_RWL<11>_XI962/MM8_g N_RBL<10>_XI962/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI962/MM7 N_XI962/NET08_XI962/MM7_d N_XI962/QB_XI962/MM7_g N_GND_XI962/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI962/MM10 N_WBL<10>_XI962/MM10_d N_WWLB<11>_XI962/MM10_g
+ N_XI962/Q_XI962/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI962/MM11 N_WBLB<10>_XI962/MM11_d N_WWLB<11>_XI962/MM11_g
+ N_XI962/QB_XI962/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI962/MM1 N_XI962/Q_XI962/MM1_d N_XI962/QB_XI962/MM1_g N_GND_XI962/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI962/MM0 N_XI962/QB_XI962/MM0_d N_XI962/Q_XI962/MM0_g N_GND_XI962/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI962/MM9 N_XI962/NET08_XI962/MM9_d N_RWLB<11>_XI962/MM9_g
+ N_RBL<10>_XI962/MM9_s N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI962/MM6 N_XI962/NET08_XI962/MM6_d N_XI962/QB_XI962/MM6_g N_VDD_XI962/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI962/MM5 N_XI962/Q_XI962/MM5_d N_XI962/QB_XI962/MM5_g N_VDD_XI962/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI962/MM4 N_XI962/QB_XI962/MM4_d N_XI962/Q_XI962/MM4_g N_VDD_XI962/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI961/MM8 N_XI961/NET08_XI961/MM8_d N_RWL<11>_XI961/MM8_g N_RBL<11>_XI961/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI961/MM7 N_XI961/NET08_XI961/MM7_d N_XI961/QB_XI961/MM7_g N_GND_XI961/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI961/MM10 N_WBL<11>_XI961/MM10_d N_WWLB<11>_XI961/MM10_g
+ N_XI961/Q_XI961/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI961/MM11 N_WBLB<11>_XI961/MM11_d N_WWLB<11>_XI961/MM11_g
+ N_XI961/QB_XI961/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI961/MM1 N_XI961/Q_XI961/MM1_d N_XI961/QB_XI961/MM1_g N_GND_XI961/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI961/MM0 N_XI961/QB_XI961/MM0_d N_XI961/Q_XI961/MM0_g N_GND_XI961/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI961/MM9 N_XI961/NET08_XI961/MM9_d N_RWLB<11>_XI961/MM9_g
+ N_RBL<11>_XI961/MM9_s N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI961/MM6 N_XI961/NET08_XI961/MM6_d N_XI961/QB_XI961/MM6_g N_VDD_XI961/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI961/MM5 N_XI961/Q_XI961/MM5_d N_XI961/QB_XI961/MM5_g N_VDD_XI961/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI961/MM4 N_XI961/QB_XI961/MM4_d N_XI961/Q_XI961/MM4_g N_VDD_XI961/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI960/MM8 N_XI960/NET08_XI960/MM8_d N_RWL<11>_XI960/MM8_g N_RBL<12>_XI960/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI960/MM7 N_XI960/NET08_XI960/MM7_d N_XI960/QB_XI960/MM7_g N_GND_XI960/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI960/MM10 N_WBL<12>_XI960/MM10_d N_WWLB<11>_XI960/MM10_g
+ N_XI960/Q_XI960/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI960/MM11 N_WBLB<12>_XI960/MM11_d N_WWLB<11>_XI960/MM11_g
+ N_XI960/QB_XI960/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI960/MM1 N_XI960/Q_XI960/MM1_d N_XI960/QB_XI960/MM1_g N_GND_XI960/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI960/MM0 N_XI960/QB_XI960/MM0_d N_XI960/Q_XI960/MM0_g N_GND_XI960/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI960/MM9 N_XI960/NET08_XI960/MM9_d N_RWLB<11>_XI960/MM9_g
+ N_RBL<12>_XI960/MM9_s N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI960/MM6 N_XI960/NET08_XI960/MM6_d N_XI960/QB_XI960/MM6_g N_VDD_XI960/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI960/MM5 N_XI960/Q_XI960/MM5_d N_XI960/QB_XI960/MM5_g N_VDD_XI960/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI960/MM4 N_XI960/QB_XI960/MM4_d N_XI960/Q_XI960/MM4_g N_VDD_XI960/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI959/MM8 N_XI959/NET08_XI959/MM8_d N_RWL<11>_XI959/MM8_g N_RBL<13>_XI959/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI959/MM7 N_XI959/NET08_XI959/MM7_d N_XI959/QB_XI959/MM7_g N_GND_XI959/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI959/MM10 N_WBL<13>_XI959/MM10_d N_WWLB<11>_XI959/MM10_g
+ N_XI959/Q_XI959/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI959/MM11 N_WBLB<13>_XI959/MM11_d N_WWLB<11>_XI959/MM11_g
+ N_XI959/QB_XI959/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI959/MM1 N_XI959/Q_XI959/MM1_d N_XI959/QB_XI959/MM1_g N_GND_XI959/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI959/MM0 N_XI959/QB_XI959/MM0_d N_XI959/Q_XI959/MM0_g N_GND_XI959/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI959/MM9 N_XI959/NET08_XI959/MM9_d N_RWLB<11>_XI959/MM9_g
+ N_RBL<13>_XI959/MM9_s N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI959/MM6 N_XI959/NET08_XI959/MM6_d N_XI959/QB_XI959/MM6_g N_VDD_XI959/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI959/MM5 N_XI959/Q_XI959/MM5_d N_XI959/QB_XI959/MM5_g N_VDD_XI959/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI959/MM4 N_XI959/QB_XI959/MM4_d N_XI959/Q_XI959/MM4_g N_VDD_XI959/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI958/MM8 N_XI958/NET08_XI958/MM8_d N_RWL<11>_XI958/MM8_g N_RBL<14>_XI958/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI958/MM7 N_XI958/NET08_XI958/MM7_d N_XI958/QB_XI958/MM7_g N_GND_XI958/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI958/MM10 N_WBL<14>_XI958/MM10_d N_WWLB<11>_XI958/MM10_g
+ N_XI958/Q_XI958/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI958/MM11 N_WBLB<14>_XI958/MM11_d N_WWLB<11>_XI958/MM11_g
+ N_XI958/QB_XI958/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI958/MM1 N_XI958/Q_XI958/MM1_d N_XI958/QB_XI958/MM1_g N_GND_XI958/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI958/MM0 N_XI958/QB_XI958/MM0_d N_XI958/Q_XI958/MM0_g N_GND_XI958/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI958/MM9 N_XI958/NET08_XI958/MM9_d N_RWLB<11>_XI958/MM9_g
+ N_RBL<14>_XI958/MM9_s N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI958/MM6 N_XI958/NET08_XI958/MM6_d N_XI958/QB_XI958/MM6_g N_VDD_XI958/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI958/MM5 N_XI958/Q_XI958/MM5_d N_XI958/QB_XI958/MM5_g N_VDD_XI958/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI958/MM4 N_XI958/QB_XI958/MM4_d N_XI958/Q_XI958/MM4_g N_VDD_XI958/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI983/MM8 N_XI983/NET08_XI983/MM8_d N_RWL<12>_XI983/MM8_g N_RBL<5>_XI983/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI983/MM7 N_XI983/NET08_XI983/MM7_d N_XI983/QB_XI983/MM7_g N_GND_XI983/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI983/MM10 N_WBL<5>_XI983/MM10_d N_WWLB<12>_XI983/MM10_g N_XI983/Q_XI983/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI983/MM11 N_WBLB<5>_XI983/MM11_d N_WWLB<12>_XI983/MM11_g
+ N_XI983/QB_XI983/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI983/MM1 N_XI983/Q_XI983/MM1_d N_XI983/QB_XI983/MM1_g N_GND_XI983/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI983/MM0 N_XI983/QB_XI983/MM0_d N_XI983/Q_XI983/MM0_g N_GND_XI983/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI983/MM9 N_XI983/NET08_XI983/MM9_d N_RWLB<12>_XI983/MM9_g N_RBL<5>_XI983/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI983/MM6 N_XI983/NET08_XI983/MM6_d N_XI983/QB_XI983/MM6_g N_VDD_XI983/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI983/MM5 N_XI983/Q_XI983/MM5_d N_XI983/QB_XI983/MM5_g N_VDD_XI983/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI983/MM4 N_XI983/QB_XI983/MM4_d N_XI983/Q_XI983/MM4_g N_VDD_XI983/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI982/MM8 N_XI982/NET08_XI982/MM8_d N_RWL<12>_XI982/MM8_g N_RBL<6>_XI982/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI982/MM7 N_XI982/NET08_XI982/MM7_d N_XI982/QB_XI982/MM7_g N_GND_XI982/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI982/MM10 N_WBL<6>_XI982/MM10_d N_WWLB<12>_XI982/MM10_g N_XI982/Q_XI982/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI982/MM11 N_WBLB<6>_XI982/MM11_d N_WWLB<12>_XI982/MM11_g
+ N_XI982/QB_XI982/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI982/MM1 N_XI982/Q_XI982/MM1_d N_XI982/QB_XI982/MM1_g N_GND_XI982/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI982/MM0 N_XI982/QB_XI982/MM0_d N_XI982/Q_XI982/MM0_g N_GND_XI982/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI982/MM9 N_XI982/NET08_XI982/MM9_d N_RWLB<12>_XI982/MM9_g N_RBL<6>_XI982/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI982/MM6 N_XI982/NET08_XI982/MM6_d N_XI982/QB_XI982/MM6_g N_VDD_XI982/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI982/MM5 N_XI982/Q_XI982/MM5_d N_XI982/QB_XI982/MM5_g N_VDD_XI982/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI982/MM4 N_XI982/QB_XI982/MM4_d N_XI982/Q_XI982/MM4_g N_VDD_XI982/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI934/MM8 N_XI934/NET08_XI934/MM8_d N_RWL<9>_XI934/MM8_g N_RBL<6>_XI934/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI934/MM7 N_XI934/NET08_XI934/MM7_d N_XI934/QB_XI934/MM7_g N_GND_XI934/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI934/MM10 N_WBL<6>_XI934/MM10_d N_WWLB<9>_XI934/MM10_g N_XI934/Q_XI934/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI934/MM11 N_WBLB<6>_XI934/MM11_d N_WWLB<9>_XI934/MM11_g
+ N_XI934/QB_XI934/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI934/MM1 N_XI934/Q_XI934/MM1_d N_XI934/QB_XI934/MM1_g N_GND_XI934/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI934/MM0 N_XI934/QB_XI934/MM0_d N_XI934/Q_XI934/MM0_g N_GND_XI934/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI934/MM9 N_XI934/NET08_XI934/MM9_d N_RWLB<9>_XI934/MM9_g N_RBL<6>_XI934/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI934/MM6 N_XI934/NET08_XI934/MM6_d N_XI934/QB_XI934/MM6_g N_VDD_XI934/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI934/MM5 N_XI934/Q_XI934/MM5_d N_XI934/QB_XI934/MM5_g N_VDD_XI934/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI934/MM4 N_XI934/QB_XI934/MM4_d N_XI934/Q_XI934/MM4_g N_VDD_XI934/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI933/MM8 N_XI933/NET08_XI933/MM8_d N_RWL<9>_XI933/MM8_g N_RBL<7>_XI933/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI933/MM7 N_XI933/NET08_XI933/MM7_d N_XI933/QB_XI933/MM7_g N_GND_XI933/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI933/MM10 N_WBL<7>_XI933/MM10_d N_WWLB<9>_XI933/MM10_g N_XI933/Q_XI933/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI933/MM11 N_WBLB<7>_XI933/MM11_d N_WWLB<9>_XI933/MM11_g
+ N_XI933/QB_XI933/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI933/MM1 N_XI933/Q_XI933/MM1_d N_XI933/QB_XI933/MM1_g N_GND_XI933/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI933/MM0 N_XI933/QB_XI933/MM0_d N_XI933/Q_XI933/MM0_g N_GND_XI933/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI933/MM9 N_XI933/NET08_XI933/MM9_d N_RWLB<9>_XI933/MM9_g N_RBL<7>_XI933/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI933/MM6 N_XI933/NET08_XI933/MM6_d N_XI933/QB_XI933/MM6_g N_VDD_XI933/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI933/MM5 N_XI933/Q_XI933/MM5_d N_XI933/QB_XI933/MM5_g N_VDD_XI933/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI933/MM4 N_XI933/QB_XI933/MM4_d N_XI933/Q_XI933/MM4_g N_VDD_XI933/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI932/MM8 N_XI932/NET08_XI932/MM8_d N_RWL<9>_XI932/MM8_g N_RBL<8>_XI932/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI932/MM7 N_XI932/NET08_XI932/MM7_d N_XI932/QB_XI932/MM7_g N_GND_XI932/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI932/MM10 N_WBL<8>_XI932/MM10_d N_WWLB<9>_XI932/MM10_g N_XI932/Q_XI932/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI932/MM11 N_WBLB<8>_XI932/MM11_d N_WWLB<9>_XI932/MM11_g
+ N_XI932/QB_XI932/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI932/MM1 N_XI932/Q_XI932/MM1_d N_XI932/QB_XI932/MM1_g N_GND_XI932/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI932/MM0 N_XI932/QB_XI932/MM0_d N_XI932/Q_XI932/MM0_g N_GND_XI932/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI932/MM9 N_XI932/NET08_XI932/MM9_d N_RWLB<9>_XI932/MM9_g N_RBL<8>_XI932/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI932/MM6 N_XI932/NET08_XI932/MM6_d N_XI932/QB_XI932/MM6_g N_VDD_XI932/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI932/MM5 N_XI932/Q_XI932/MM5_d N_XI932/QB_XI932/MM5_g N_VDD_XI932/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI932/MM4 N_XI932/QB_XI932/MM4_d N_XI932/Q_XI932/MM4_g N_VDD_XI932/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI935/MM8 N_XI935/NET08_XI935/MM8_d N_RWL<9>_XI935/MM8_g N_RBL<5>_XI935/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI935/MM7 N_XI935/NET08_XI935/MM7_d N_XI935/QB_XI935/MM7_g N_GND_XI935/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI935/MM10 N_WBL<5>_XI935/MM10_d N_WWLB<9>_XI935/MM10_g N_XI935/Q_XI935/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI935/MM11 N_WBLB<5>_XI935/MM11_d N_WWLB<9>_XI935/MM11_g
+ N_XI935/QB_XI935/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI935/MM1 N_XI935/Q_XI935/MM1_d N_XI935/QB_XI935/MM1_g N_GND_XI935/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI935/MM0 N_XI935/QB_XI935/MM0_d N_XI935/Q_XI935/MM0_g N_GND_XI935/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI935/MM9 N_XI935/NET08_XI935/MM9_d N_RWLB<9>_XI935/MM9_g N_RBL<5>_XI935/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI935/MM6 N_XI935/NET08_XI935/MM6_d N_XI935/QB_XI935/MM6_g N_VDD_XI935/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI935/MM5 N_XI935/Q_XI935/MM5_d N_XI935/QB_XI935/MM5_g N_VDD_XI935/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI935/MM4 N_XI935/QB_XI935/MM4_d N_XI935/Q_XI935/MM4_g N_VDD_XI935/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1032/MM8 N_XI1032/NET08_XI1032/MM8_d N_RWL<15>_XI1032/MM8_g
+ N_RBL<4>_XI1032/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1032/MM7 N_XI1032/NET08_XI1032/MM7_d N_XI1032/QB_XI1032/MM7_g
+ N_GND_XI1032/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1032/MM10 N_WBL<4>_XI1032/MM10_d N_WWLB<15>_XI1032/MM10_g
+ N_XI1032/Q_XI1032/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1032/MM11 N_WBLB<4>_XI1032/MM11_d N_WWLB<15>_XI1032/MM11_g
+ N_XI1032/QB_XI1032/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1032/MM1 N_XI1032/Q_XI1032/MM1_d N_XI1032/QB_XI1032/MM1_g N_GND_XI1032/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1032/MM0 N_XI1032/QB_XI1032/MM0_d N_XI1032/Q_XI1032/MM0_g N_GND_XI1032/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1032/MM9 N_XI1032/NET08_XI1032/MM9_d N_RWLB<15>_XI1032/MM9_g
+ N_RBL<4>_XI1032/MM9_s N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1032/MM6 N_XI1032/NET08_XI1032/MM6_d N_XI1032/QB_XI1032/MM6_g
+ N_VDD_XI1032/MM6_s N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1032/MM5 N_XI1032/Q_XI1032/MM5_d N_XI1032/QB_XI1032/MM5_g N_VDD_XI1032/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1032/MM4 N_XI1032/QB_XI1032/MM4_d N_XI1032/Q_XI1032/MM4_g N_VDD_XI1032/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI995/MM8 N_XI995/NET08_XI995/MM8_d N_RWL<13>_XI995/MM8_g N_RBL<9>_XI995/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI995/MM7 N_XI995/NET08_XI995/MM7_d N_XI995/QB_XI995/MM7_g N_GND_XI995/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI995/MM10 N_WBL<9>_XI995/MM10_d N_WWLB<13>_XI995/MM10_g N_XI995/Q_XI995/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI995/MM11 N_WBLB<9>_XI995/MM11_d N_WWLB<13>_XI995/MM11_g
+ N_XI995/QB_XI995/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI995/MM1 N_XI995/Q_XI995/MM1_d N_XI995/QB_XI995/MM1_g N_GND_XI995/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI995/MM0 N_XI995/QB_XI995/MM0_d N_XI995/Q_XI995/MM0_g N_GND_XI995/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI995/MM9 N_XI995/NET08_XI995/MM9_d N_RWLB<13>_XI995/MM9_g N_RBL<9>_XI995/MM9_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI995/MM6 N_XI995/NET08_XI995/MM6_d N_XI995/QB_XI995/MM6_g N_VDD_XI995/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI995/MM5 N_XI995/Q_XI995/MM5_d N_XI995/QB_XI995/MM5_g N_VDD_XI995/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI995/MM4 N_XI995/QB_XI995/MM4_d N_XI995/Q_XI995/MM4_g N_VDD_XI995/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI938/MM8 N_XI938/NET08_XI938/MM8_d N_RWL<9>_XI938/MM8_g N_RBL<2>_XI938/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI938/MM7 N_XI938/NET08_XI938/MM7_d N_XI938/QB_XI938/MM7_g N_GND_XI938/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI938/MM10 N_WBL<2>_XI938/MM10_d N_WWLB<9>_XI938/MM10_g N_XI938/Q_XI938/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI938/MM11 N_WBLB<2>_XI938/MM11_d N_WWLB<9>_XI938/MM11_g
+ N_XI938/QB_XI938/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI938/MM1 N_XI938/Q_XI938/MM1_d N_XI938/QB_XI938/MM1_g N_GND_XI938/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI938/MM0 N_XI938/QB_XI938/MM0_d N_XI938/Q_XI938/MM0_g N_GND_XI938/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI938/MM9 N_XI938/NET08_XI938/MM9_d N_RWLB<9>_XI938/MM9_g N_RBL<2>_XI938/MM9_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI938/MM6 N_XI938/NET08_XI938/MM6_d N_XI938/QB_XI938/MM6_g N_VDD_XI938/MM6_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI938/MM5 N_XI938/Q_XI938/MM5_d N_XI938/QB_XI938/MM5_g N_VDD_XI938/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI938/MM4 N_XI938/QB_XI938/MM4_d N_XI938/Q_XI938/MM4_g N_VDD_XI938/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI937/MM8 N_XI937/NET08_XI937/MM8_d N_RWL<9>_XI937/MM8_g N_RBL<3>_XI937/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI937/MM7 N_XI937/NET08_XI937/MM7_d N_XI937/QB_XI937/MM7_g N_GND_XI937/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI937/MM10 N_WBL<3>_XI937/MM10_d N_WWLB<9>_XI937/MM10_g N_XI937/Q_XI937/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI937/MM11 N_WBLB<3>_XI937/MM11_d N_WWLB<9>_XI937/MM11_g
+ N_XI937/QB_XI937/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI937/MM1 N_XI937/Q_XI937/MM1_d N_XI937/QB_XI937/MM1_g N_GND_XI937/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI937/MM0 N_XI937/QB_XI937/MM0_d N_XI937/Q_XI937/MM0_g N_GND_XI937/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI937/MM9 N_XI937/NET08_XI937/MM9_d N_RWLB<9>_XI937/MM9_g N_RBL<3>_XI937/MM9_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI937/MM6 N_XI937/NET08_XI937/MM6_d N_XI937/QB_XI937/MM6_g N_VDD_XI937/MM6_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI937/MM5 N_XI937/Q_XI937/MM5_d N_XI937/QB_XI937/MM5_g N_VDD_XI937/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI937/MM4 N_XI937/QB_XI937/MM4_d N_XI937/Q_XI937/MM4_g N_VDD_XI937/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI936/MM8 N_XI936/NET08_XI936/MM8_d N_RWL<9>_XI936/MM8_g N_RBL<4>_XI936/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI936/MM7 N_XI936/NET08_XI936/MM7_d N_XI936/QB_XI936/MM7_g N_GND_XI936/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI936/MM10 N_WBL<4>_XI936/MM10_d N_WWLB<9>_XI936/MM10_g N_XI936/Q_XI936/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI936/MM11 N_WBLB<4>_XI936/MM11_d N_WWLB<9>_XI936/MM11_g
+ N_XI936/QB_XI936/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI936/MM1 N_XI936/Q_XI936/MM1_d N_XI936/QB_XI936/MM1_g N_GND_XI936/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI936/MM0 N_XI936/QB_XI936/MM0_d N_XI936/Q_XI936/MM0_g N_GND_XI936/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI936/MM9 N_XI936/NET08_XI936/MM9_d N_RWLB<9>_XI936/MM9_g N_RBL<4>_XI936/MM9_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI936/MM6 N_XI936/NET08_XI936/MM6_d N_XI936/QB_XI936/MM6_g N_VDD_XI936/MM6_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI936/MM5 N_XI936/Q_XI936/MM5_d N_XI936/QB_XI936/MM5_g N_VDD_XI936/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI936/MM4 N_XI936/QB_XI936/MM4_d N_XI936/Q_XI936/MM4_g N_VDD_XI936/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI939/MM8 N_XI939/NET08_XI939/MM8_d N_RWL<9>_XI939/MM8_g N_RBL<1>_XI939/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI939/MM7 N_XI939/NET08_XI939/MM7_d N_XI939/QB_XI939/MM7_g N_GND_XI939/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI939/MM10 N_WBL<1>_XI939/MM10_d N_WWLB<9>_XI939/MM10_g N_XI939/Q_XI939/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI939/MM11 N_WBLB<1>_XI939/MM11_d N_WWLB<9>_XI939/MM11_g
+ N_XI939/QB_XI939/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI939/MM1 N_XI939/Q_XI939/MM1_d N_XI939/QB_XI939/MM1_g N_GND_XI939/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI939/MM0 N_XI939/QB_XI939/MM0_d N_XI939/Q_XI939/MM0_g N_GND_XI939/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI939/MM9 N_XI939/NET08_XI939/MM9_d N_RWLB<9>_XI939/MM9_g N_RBL<1>_XI939/MM9_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI939/MM6 N_XI939/NET08_XI939/MM6_d N_XI939/QB_XI939/MM6_g N_VDD_XI939/MM6_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI939/MM5 N_XI939/Q_XI939/MM5_d N_XI939/QB_XI939/MM5_g N_VDD_XI939/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI939/MM4 N_XI939/QB_XI939/MM4_d N_XI939/Q_XI939/MM4_g N_VDD_XI939/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI956/MM8 N_XI956/NET08_XI956/MM8_d N_RWL<10>_XI956/MM8_g N_RBL<0>_XI956/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI956/MM7 N_XI956/NET08_XI956/MM7_d N_XI956/QB_XI956/MM7_g N_GND_XI956/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI956/MM10 N_WBL<0>_XI956/MM10_d N_WWLB<10>_XI956/MM10_g N_XI956/Q_XI956/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI956/MM11 N_WBLB<0>_XI956/MM11_d N_WWLB<10>_XI956/MM11_g
+ N_XI956/QB_XI956/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI956/MM1 N_XI956/Q_XI956/MM1_d N_XI956/QB_XI956/MM1_g N_GND_XI956/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI956/MM0 N_XI956/QB_XI956/MM0_d N_XI956/Q_XI956/MM0_g N_GND_XI956/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI956/MM9 N_XI956/NET08_XI956/MM9_d N_RWLB<10>_XI956/MM9_g N_RBL<0>_XI956/MM9_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI956/MM6 N_XI956/NET08_XI956/MM6_d N_XI956/QB_XI956/MM6_g N_VDD_XI956/MM6_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI956/MM5 N_XI956/Q_XI956/MM5_d N_XI956/QB_XI956/MM5_g N_VDD_XI956/MM5_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI956/MM4 N_XI956/QB_XI956/MM4_d N_XI956/Q_XI956/MM4_g N_VDD_XI956/MM4_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI955/MM8 N_XI955/NET08_XI955/MM8_d N_RWL<10>_XI955/MM8_g N_RBL<1>_XI955/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI955/MM7 N_XI955/NET08_XI955/MM7_d N_XI955/QB_XI955/MM7_g N_GND_XI955/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI955/MM10 N_WBL<1>_XI955/MM10_d N_WWLB<10>_XI955/MM10_g N_XI955/Q_XI955/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI955/MM11 N_WBLB<1>_XI955/MM11_d N_WWLB<10>_XI955/MM11_g
+ N_XI955/QB_XI955/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI955/MM1 N_XI955/Q_XI955/MM1_d N_XI955/QB_XI955/MM1_g N_GND_XI955/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI955/MM0 N_XI955/QB_XI955/MM0_d N_XI955/Q_XI955/MM0_g N_GND_XI955/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI955/MM9 N_XI955/NET08_XI955/MM9_d N_RWLB<10>_XI955/MM9_g N_RBL<1>_XI955/MM9_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI955/MM6 N_XI955/NET08_XI955/MM6_d N_XI955/QB_XI955/MM6_g N_VDD_XI955/MM6_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI955/MM5 N_XI955/Q_XI955/MM5_d N_XI955/QB_XI955/MM5_g N_VDD_XI955/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI955/MM4 N_XI955/QB_XI955/MM4_d N_XI955/Q_XI955/MM4_g N_VDD_XI955/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI954/MM8 N_XI954/NET08_XI954/MM8_d N_RWL<10>_XI954/MM8_g N_RBL<2>_XI954/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI954/MM7 N_XI954/NET08_XI954/MM7_d N_XI954/QB_XI954/MM7_g N_GND_XI954/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI954/MM10 N_WBL<2>_XI954/MM10_d N_WWLB<10>_XI954/MM10_g N_XI954/Q_XI954/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI954/MM11 N_WBLB<2>_XI954/MM11_d N_WWLB<10>_XI954/MM11_g
+ N_XI954/QB_XI954/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI954/MM1 N_XI954/Q_XI954/MM1_d N_XI954/QB_XI954/MM1_g N_GND_XI954/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI954/MM0 N_XI954/QB_XI954/MM0_d N_XI954/Q_XI954/MM0_g N_GND_XI954/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI954/MM9 N_XI954/NET08_XI954/MM9_d N_RWLB<10>_XI954/MM9_g N_RBL<2>_XI954/MM9_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI954/MM6 N_XI954/NET08_XI954/MM6_d N_XI954/QB_XI954/MM6_g N_VDD_XI954/MM6_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI954/MM5 N_XI954/Q_XI954/MM5_d N_XI954/QB_XI954/MM5_g N_VDD_XI954/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI954/MM4 N_XI954/QB_XI954/MM4_d N_XI954/Q_XI954/MM4_g N_VDD_XI954/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI953/MM8 N_XI953/NET08_XI953/MM8_d N_RWL<10>_XI953/MM8_g N_RBL<3>_XI953/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI953/MM7 N_XI953/NET08_XI953/MM7_d N_XI953/QB_XI953/MM7_g N_GND_XI953/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI953/MM10 N_WBL<3>_XI953/MM10_d N_WWLB<10>_XI953/MM10_g N_XI953/Q_XI953/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI953/MM11 N_WBLB<3>_XI953/MM11_d N_WWLB<10>_XI953/MM11_g
+ N_XI953/QB_XI953/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI953/MM1 N_XI953/Q_XI953/MM1_d N_XI953/QB_XI953/MM1_g N_GND_XI953/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI953/MM0 N_XI953/QB_XI953/MM0_d N_XI953/Q_XI953/MM0_g N_GND_XI953/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI953/MM9 N_XI953/NET08_XI953/MM9_d N_RWLB<10>_XI953/MM9_g N_RBL<3>_XI953/MM9_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI953/MM6 N_XI953/NET08_XI953/MM6_d N_XI953/QB_XI953/MM6_g N_VDD_XI953/MM6_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI953/MM5 N_XI953/Q_XI953/MM5_d N_XI953/QB_XI953/MM5_g N_VDD_XI953/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI953/MM4 N_XI953/QB_XI953/MM4_d N_XI953/Q_XI953/MM4_g N_VDD_XI953/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI952/MM8 N_XI952/NET08_XI952/MM8_d N_RWL<10>_XI952/MM8_g N_RBL<4>_XI952/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI952/MM7 N_XI952/NET08_XI952/MM7_d N_XI952/QB_XI952/MM7_g N_GND_XI952/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI952/MM10 N_WBL<4>_XI952/MM10_d N_WWLB<10>_XI952/MM10_g N_XI952/Q_XI952/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI952/MM11 N_WBLB<4>_XI952/MM11_d N_WWLB<10>_XI952/MM11_g
+ N_XI952/QB_XI952/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI952/MM1 N_XI952/Q_XI952/MM1_d N_XI952/QB_XI952/MM1_g N_GND_XI952/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI952/MM0 N_XI952/QB_XI952/MM0_d N_XI952/Q_XI952/MM0_g N_GND_XI952/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI952/MM9 N_XI952/NET08_XI952/MM9_d N_RWLB<10>_XI952/MM9_g N_RBL<4>_XI952/MM9_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI952/MM6 N_XI952/NET08_XI952/MM6_d N_XI952/QB_XI952/MM6_g N_VDD_XI952/MM6_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI952/MM5 N_XI952/Q_XI952/MM5_d N_XI952/QB_XI952/MM5_g N_VDD_XI952/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI952/MM4 N_XI952/QB_XI952/MM4_d N_XI952/Q_XI952/MM4_g N_VDD_XI952/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI957/MM8 N_XI957/NET08_XI957/MM8_d N_RWL<10>_XI957/MM8_g N_RBL<15>_XI957/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI957/MM7 N_XI957/NET08_XI957/MM7_d N_XI957/QB_XI957/MM7_g N_GND_XI957/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI957/MM10 N_WBL<15>_XI957/MM10_d N_WWLB<10>_XI957/MM10_g
+ N_XI957/Q_XI957/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI957/MM11 N_WBLB<15>_XI957/MM11_d N_WWLB<10>_XI957/MM11_g
+ N_XI957/QB_XI957/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI957/MM1 N_XI957/Q_XI957/MM1_d N_XI957/QB_XI957/MM1_g N_GND_XI957/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI957/MM0 N_XI957/QB_XI957/MM0_d N_XI957/Q_XI957/MM0_g N_GND_XI957/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI957/MM9 N_XI957/NET08_XI957/MM9_d N_RWLB<10>_XI957/MM9_g
+ N_RBL<15>_XI957/MM9_s N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI957/MM6 N_XI957/NET08_XI957/MM6_d N_XI957/QB_XI957/MM6_g N_VDD_XI957/MM6_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI957/MM5 N_XI957/Q_XI957/MM5_d N_XI957/QB_XI957/MM5_g N_VDD_XI957/MM5_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI957/MM4 N_XI957/QB_XI957/MM4_d N_XI957/Q_XI957/MM4_g N_VDD_XI957/MM4_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI979/MM8 N_XI979/NET08_XI979/MM8_d N_RWL<12>_XI979/MM8_g N_RBL<9>_XI979/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI979/MM7 N_XI979/NET08_XI979/MM7_d N_XI979/QB_XI979/MM7_g N_GND_XI979/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI979/MM10 N_WBL<9>_XI979/MM10_d N_WWLB<12>_XI979/MM10_g N_XI979/Q_XI979/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI979/MM11 N_WBLB<9>_XI979/MM11_d N_WWLB<12>_XI979/MM11_g
+ N_XI979/QB_XI979/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI979/MM1 N_XI979/Q_XI979/MM1_d N_XI979/QB_XI979/MM1_g N_GND_XI979/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI979/MM0 N_XI979/QB_XI979/MM0_d N_XI979/Q_XI979/MM0_g N_GND_XI979/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI979/MM9 N_XI979/NET08_XI979/MM9_d N_RWLB<12>_XI979/MM9_g N_RBL<9>_XI979/MM9_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI979/MM6 N_XI979/NET08_XI979/MM6_d N_XI979/QB_XI979/MM6_g N_VDD_XI979/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI979/MM5 N_XI979/Q_XI979/MM5_d N_XI979/QB_XI979/MM5_g N_VDD_XI979/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI979/MM4 N_XI979/QB_XI979/MM4_d N_XI979/Q_XI979/MM4_g N_VDD_XI979/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI900/MM8 N_XI900/NET08_XI900/MM8_d N_RWL<7>_XI900/MM8_g N_RBL<8>_XI900/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI900/MM7 N_XI900/NET08_XI900/MM7_d N_XI900/QB_XI900/MM7_g N_GND_XI900/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI900/MM10 N_WBL<8>_XI900/MM10_d N_WWLB<7>_XI900/MM10_g N_XI900/Q_XI900/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI900/MM11 N_WBLB<8>_XI900/MM11_d N_WWLB<7>_XI900/MM11_g
+ N_XI900/QB_XI900/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI900/MM1 N_XI900/Q_XI900/MM1_d N_XI900/QB_XI900/MM1_g N_GND_XI900/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI900/MM0 N_XI900/QB_XI900/MM0_d N_XI900/Q_XI900/MM0_g N_GND_XI900/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI900/MM9 N_XI900/NET08_XI900/MM9_d N_RWLB<7>_XI900/MM9_g N_RBL<8>_XI900/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI900/MM6 N_XI900/NET08_XI900/MM6_d N_XI900/QB_XI900/MM6_g N_VDD_XI900/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI900/MM5 N_XI900/Q_XI900/MM5_d N_XI900/QB_XI900/MM5_g N_VDD_XI900/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI900/MM4 N_XI900/QB_XI900/MM4_d N_XI900/Q_XI900/MM4_g N_VDD_XI900/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI931/MM8 N_XI931/NET08_XI931/MM8_d N_RWL<9>_XI931/MM8_g N_RBL<9>_XI931/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI931/MM7 N_XI931/NET08_XI931/MM7_d N_XI931/QB_XI931/MM7_g N_GND_XI931/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI931/MM10 N_WBL<9>_XI931/MM10_d N_WWLB<9>_XI931/MM10_g N_XI931/Q_XI931/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI931/MM11 N_WBLB<9>_XI931/MM11_d N_WWLB<9>_XI931/MM11_g
+ N_XI931/QB_XI931/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI931/MM1 N_XI931/Q_XI931/MM1_d N_XI931/QB_XI931/MM1_g N_GND_XI931/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI931/MM0 N_XI931/QB_XI931/MM0_d N_XI931/Q_XI931/MM0_g N_GND_XI931/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI931/MM9 N_XI931/NET08_XI931/MM9_d N_RWLB<9>_XI931/MM9_g N_RBL<9>_XI931/MM9_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI931/MM6 N_XI931/NET08_XI931/MM6_d N_XI931/QB_XI931/MM6_g N_VDD_XI931/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI931/MM5 N_XI931/Q_XI931/MM5_d N_XI931/QB_XI931/MM5_g N_VDD_XI931/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI931/MM4 N_XI931/QB_XI931/MM4_d N_XI931/Q_XI931/MM4_g N_VDD_XI931/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI930/MM8 N_XI930/NET08_XI930/MM8_d N_RWL<9>_XI930/MM8_g N_RBL<10>_XI930/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI930/MM7 N_XI930/NET08_XI930/MM7_d N_XI930/QB_XI930/MM7_g N_GND_XI930/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI930/MM10 N_WBL<10>_XI930/MM10_d N_WWLB<9>_XI930/MM10_g N_XI930/Q_XI930/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI930/MM11 N_WBLB<10>_XI930/MM11_d N_WWLB<9>_XI930/MM11_g
+ N_XI930/QB_XI930/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI930/MM1 N_XI930/Q_XI930/MM1_d N_XI930/QB_XI930/MM1_g N_GND_XI930/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI930/MM0 N_XI930/QB_XI930/MM0_d N_XI930/Q_XI930/MM0_g N_GND_XI930/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI930/MM9 N_XI930/NET08_XI930/MM9_d N_RWLB<9>_XI930/MM9_g N_RBL<10>_XI930/MM9_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI930/MM6 N_XI930/NET08_XI930/MM6_d N_XI930/QB_XI930/MM6_g N_VDD_XI930/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI930/MM5 N_XI930/Q_XI930/MM5_d N_XI930/QB_XI930/MM5_g N_VDD_XI930/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI930/MM4 N_XI930/QB_XI930/MM4_d N_XI930/Q_XI930/MM4_g N_VDD_XI930/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI929/MM8 N_XI929/NET08_XI929/MM8_d N_RWL<9>_XI929/MM8_g N_RBL<11>_XI929/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI929/MM7 N_XI929/NET08_XI929/MM7_d N_XI929/QB_XI929/MM7_g N_GND_XI929/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI929/MM10 N_WBL<11>_XI929/MM10_d N_WWLB<9>_XI929/MM10_g N_XI929/Q_XI929/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI929/MM11 N_WBLB<11>_XI929/MM11_d N_WWLB<9>_XI929/MM11_g
+ N_XI929/QB_XI929/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI929/MM1 N_XI929/Q_XI929/MM1_d N_XI929/QB_XI929/MM1_g N_GND_XI929/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI929/MM0 N_XI929/QB_XI929/MM0_d N_XI929/Q_XI929/MM0_g N_GND_XI929/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI929/MM9 N_XI929/NET08_XI929/MM9_d N_RWLB<9>_XI929/MM9_g N_RBL<11>_XI929/MM9_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI929/MM6 N_XI929/NET08_XI929/MM6_d N_XI929/QB_XI929/MM6_g N_VDD_XI929/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI929/MM5 N_XI929/Q_XI929/MM5_d N_XI929/QB_XI929/MM5_g N_VDD_XI929/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI929/MM4 N_XI929/QB_XI929/MM4_d N_XI929/Q_XI929/MM4_g N_VDD_XI929/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI928/MM8 N_XI928/NET08_XI928/MM8_d N_RWL<9>_XI928/MM8_g N_RBL<12>_XI928/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI928/MM7 N_XI928/NET08_XI928/MM7_d N_XI928/QB_XI928/MM7_g N_GND_XI928/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI928/MM10 N_WBL<12>_XI928/MM10_d N_WWLB<9>_XI928/MM10_g N_XI928/Q_XI928/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI928/MM11 N_WBLB<12>_XI928/MM11_d N_WWLB<9>_XI928/MM11_g
+ N_XI928/QB_XI928/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI928/MM1 N_XI928/Q_XI928/MM1_d N_XI928/QB_XI928/MM1_g N_GND_XI928/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI928/MM0 N_XI928/QB_XI928/MM0_d N_XI928/Q_XI928/MM0_g N_GND_XI928/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI928/MM9 N_XI928/NET08_XI928/MM9_d N_RWLB<9>_XI928/MM9_g N_RBL<12>_XI928/MM9_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI928/MM6 N_XI928/NET08_XI928/MM6_d N_XI928/QB_XI928/MM6_g N_VDD_XI928/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI928/MM5 N_XI928/Q_XI928/MM5_d N_XI928/QB_XI928/MM5_g N_VDD_XI928/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI928/MM4 N_XI928/QB_XI928/MM4_d N_XI928/Q_XI928/MM4_g N_VDD_XI928/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1031/MM8 N_XI1031/NET08_XI1031/MM8_d N_RWL<15>_XI1031/MM8_g
+ N_RBL<5>_XI1031/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1031/MM7 N_XI1031/NET08_XI1031/MM7_d N_XI1031/QB_XI1031/MM7_g
+ N_GND_XI1031/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1031/MM10 N_WBL<5>_XI1031/MM10_d N_WWLB<15>_XI1031/MM10_g
+ N_XI1031/Q_XI1031/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1031/MM11 N_WBLB<5>_XI1031/MM11_d N_WWLB<15>_XI1031/MM11_g
+ N_XI1031/QB_XI1031/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1031/MM1 N_XI1031/Q_XI1031/MM1_d N_XI1031/QB_XI1031/MM1_g N_GND_XI1031/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1031/MM0 N_XI1031/QB_XI1031/MM0_d N_XI1031/Q_XI1031/MM0_g N_GND_XI1031/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1031/MM9 N_XI1031/NET08_XI1031/MM9_d N_RWLB<15>_XI1031/MM9_g
+ N_RBL<5>_XI1031/MM9_s N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1031/MM6 N_XI1031/NET08_XI1031/MM6_d N_XI1031/QB_XI1031/MM6_g
+ N_VDD_XI1031/MM6_s N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1031/MM5 N_XI1031/Q_XI1031/MM5_d N_XI1031/QB_XI1031/MM5_g N_VDD_XI1031/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1031/MM4 N_XI1031/QB_XI1031/MM4_d N_XI1031/Q_XI1031/MM4_g N_VDD_XI1031/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI996/MM8 N_XI996/NET08_XI996/MM8_d N_RWL<13>_XI996/MM8_g N_RBL<8>_XI996/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI996/MM7 N_XI996/NET08_XI996/MM7_d N_XI996/QB_XI996/MM7_g N_GND_XI996/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI996/MM10 N_WBL<8>_XI996/MM10_d N_WWLB<13>_XI996/MM10_g N_XI996/Q_XI996/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI996/MM11 N_WBLB<8>_XI996/MM11_d N_WWLB<13>_XI996/MM11_g
+ N_XI996/QB_XI996/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI996/MM1 N_XI996/Q_XI996/MM1_d N_XI996/QB_XI996/MM1_g N_GND_XI996/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI996/MM0 N_XI996/QB_XI996/MM0_d N_XI996/Q_XI996/MM0_g N_GND_XI996/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI996/MM9 N_XI996/NET08_XI996/MM9_d N_RWLB<13>_XI996/MM9_g N_RBL<8>_XI996/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI996/MM6 N_XI996/NET08_XI996/MM6_d N_XI996/QB_XI996/MM6_g N_VDD_XI996/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI996/MM5 N_XI996/Q_XI996/MM5_d N_XI996/QB_XI996/MM5_g N_VDD_XI996/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI996/MM4 N_XI996/QB_XI996/MM4_d N_XI996/Q_XI996/MM4_g N_VDD_XI996/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI875/MM8 N_XI875/NET08_XI875/MM8_d N_RWL<5>_XI875/MM8_g N_RBL<1>_XI875/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI875/MM7 N_XI875/NET08_XI875/MM7_d N_XI875/QB_XI875/MM7_g N_GND_XI875/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI875/MM10 N_WBL<1>_XI875/MM10_d N_WWLB<5>_XI875/MM10_g N_XI875/Q_XI875/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI875/MM11 N_WBLB<1>_XI875/MM11_d N_WWLB<5>_XI875/MM11_g
+ N_XI875/QB_XI875/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI875/MM1 N_XI875/Q_XI875/MM1_d N_XI875/QB_XI875/MM1_g N_GND_XI875/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI875/MM0 N_XI875/QB_XI875/MM0_d N_XI875/Q_XI875/MM0_g N_GND_XI875/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI875/MM9 N_XI875/NET08_XI875/MM9_d N_RWLB<5>_XI875/MM9_g N_RBL<1>_XI875/MM9_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI875/MM6 N_XI875/NET08_XI875/MM6_d N_XI875/QB_XI875/MM6_g N_VDD_XI875/MM6_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI875/MM5 N_XI875/Q_XI875/MM5_d N_XI875/QB_XI875/MM5_g N_VDD_XI875/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI875/MM4 N_XI875/QB_XI875/MM4_d N_XI875/Q_XI875/MM4_g N_VDD_XI875/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI874/MM8 N_XI874/NET08_XI874/MM8_d N_RWL<5>_XI874/MM8_g N_RBL<2>_XI874/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI874/MM7 N_XI874/NET08_XI874/MM7_d N_XI874/QB_XI874/MM7_g N_GND_XI874/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI874/MM10 N_WBL<2>_XI874/MM10_d N_WWLB<5>_XI874/MM10_g N_XI874/Q_XI874/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI874/MM11 N_WBLB<2>_XI874/MM11_d N_WWLB<5>_XI874/MM11_g
+ N_XI874/QB_XI874/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI874/MM1 N_XI874/Q_XI874/MM1_d N_XI874/QB_XI874/MM1_g N_GND_XI874/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI874/MM0 N_XI874/QB_XI874/MM0_d N_XI874/Q_XI874/MM0_g N_GND_XI874/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI874/MM9 N_XI874/NET08_XI874/MM9_d N_RWLB<5>_XI874/MM9_g N_RBL<2>_XI874/MM9_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI874/MM6 N_XI874/NET08_XI874/MM6_d N_XI874/QB_XI874/MM6_g N_VDD_XI874/MM6_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI874/MM5 N_XI874/Q_XI874/MM5_d N_XI874/QB_XI874/MM5_g N_VDD_XI874/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI874/MM4 N_XI874/QB_XI874/MM4_d N_XI874/Q_XI874/MM4_g N_VDD_XI874/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI873/MM8 N_XI873/NET08_XI873/MM8_d N_RWL<5>_XI873/MM8_g N_RBL<3>_XI873/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI873/MM7 N_XI873/NET08_XI873/MM7_d N_XI873/QB_XI873/MM7_g N_GND_XI873/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI873/MM10 N_WBL<3>_XI873/MM10_d N_WWLB<5>_XI873/MM10_g N_XI873/Q_XI873/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI873/MM11 N_WBLB<3>_XI873/MM11_d N_WWLB<5>_XI873/MM11_g
+ N_XI873/QB_XI873/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI873/MM1 N_XI873/Q_XI873/MM1_d N_XI873/QB_XI873/MM1_g N_GND_XI873/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI873/MM0 N_XI873/QB_XI873/MM0_d N_XI873/Q_XI873/MM0_g N_GND_XI873/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI873/MM9 N_XI873/NET08_XI873/MM9_d N_RWLB<5>_XI873/MM9_g N_RBL<3>_XI873/MM9_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI873/MM6 N_XI873/NET08_XI873/MM6_d N_XI873/QB_XI873/MM6_g N_VDD_XI873/MM6_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI873/MM5 N_XI873/Q_XI873/MM5_d N_XI873/QB_XI873/MM5_g N_VDD_XI873/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI873/MM4 N_XI873/QB_XI873/MM4_d N_XI873/Q_XI873/MM4_g N_VDD_XI873/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI872/MM8 N_XI872/NET08_XI872/MM8_d N_RWL<5>_XI872/MM8_g N_RBL<4>_XI872/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI872/MM7 N_XI872/NET08_XI872/MM7_d N_XI872/QB_XI872/MM7_g N_GND_XI872/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI872/MM10 N_WBL<4>_XI872/MM10_d N_WWLB<5>_XI872/MM10_g N_XI872/Q_XI872/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI872/MM11 N_WBLB<4>_XI872/MM11_d N_WWLB<5>_XI872/MM11_g
+ N_XI872/QB_XI872/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI872/MM1 N_XI872/Q_XI872/MM1_d N_XI872/QB_XI872/MM1_g N_GND_XI872/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI872/MM0 N_XI872/QB_XI872/MM0_d N_XI872/Q_XI872/MM0_g N_GND_XI872/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI872/MM9 N_XI872/NET08_XI872/MM9_d N_RWLB<5>_XI872/MM9_g N_RBL<4>_XI872/MM9_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI872/MM6 N_XI872/NET08_XI872/MM6_d N_XI872/QB_XI872/MM6_g N_VDD_XI872/MM6_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI872/MM5 N_XI872/Q_XI872/MM5_d N_XI872/QB_XI872/MM5_g N_VDD_XI872/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI872/MM4 N_XI872/QB_XI872/MM4_d N_XI872/Q_XI872/MM4_g N_VDD_XI872/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI911/MM8 N_XI911/NET08_XI911/MM8_d N_RWL<8>_XI911/MM8_g N_RBL<13>_XI911/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI911/MM7 N_XI911/NET08_XI911/MM7_d N_XI911/QB_XI911/MM7_g N_GND_XI911/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI911/MM10 N_WBL<13>_XI911/MM10_d N_WWLB<8>_XI911/MM10_g N_XI911/Q_XI911/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI911/MM11 N_WBLB<13>_XI911/MM11_d N_WWLB<8>_XI911/MM11_g
+ N_XI911/QB_XI911/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI911/MM1 N_XI911/Q_XI911/MM1_d N_XI911/QB_XI911/MM1_g N_GND_XI911/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI911/MM0 N_XI911/QB_XI911/MM0_d N_XI911/Q_XI911/MM0_g N_GND_XI911/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI911/MM9 N_XI911/NET08_XI911/MM9_d N_RWLB<8>_XI911/MM9_g N_RBL<13>_XI911/MM9_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI911/MM6 N_XI911/NET08_XI911/MM6_d N_XI911/QB_XI911/MM6_g N_VDD_XI911/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI911/MM5 N_XI911/Q_XI911/MM5_d N_XI911/QB_XI911/MM5_g N_VDD_XI911/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI911/MM4 N_XI911/QB_XI911/MM4_d N_XI911/Q_XI911/MM4_g N_VDD_XI911/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI910/MM8 N_XI910/NET08_XI910/MM8_d N_RWL<8>_XI910/MM8_g N_RBL<14>_XI910/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI910/MM7 N_XI910/NET08_XI910/MM7_d N_XI910/QB_XI910/MM7_g N_GND_XI910/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI910/MM10 N_WBL<14>_XI910/MM10_d N_WWLB<8>_XI910/MM10_g N_XI910/Q_XI910/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI910/MM11 N_WBLB<14>_XI910/MM11_d N_WWLB<8>_XI910/MM11_g
+ N_XI910/QB_XI910/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI910/MM1 N_XI910/Q_XI910/MM1_d N_XI910/QB_XI910/MM1_g N_GND_XI910/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI910/MM0 N_XI910/QB_XI910/MM0_d N_XI910/Q_XI910/MM0_g N_GND_XI910/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI910/MM9 N_XI910/NET08_XI910/MM9_d N_RWLB<8>_XI910/MM9_g N_RBL<14>_XI910/MM9_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI910/MM6 N_XI910/NET08_XI910/MM6_d N_XI910/QB_XI910/MM6_g N_VDD_XI910/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI910/MM5 N_XI910/Q_XI910/MM5_d N_XI910/QB_XI910/MM5_g N_VDD_XI910/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI910/MM4 N_XI910/QB_XI910/MM4_d N_XI910/Q_XI910/MM4_g N_VDD_XI910/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI909/MM8 N_XI909/NET08_XI909/MM8_d N_RWL<7>_XI909/MM8_g N_RBL<15>_XI909/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI909/MM7 N_XI909/NET08_XI909/MM7_d N_XI909/QB_XI909/MM7_g N_GND_XI909/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI909/MM10 N_WBL<15>_XI909/MM10_d N_WWLB<7>_XI909/MM10_g N_XI909/Q_XI909/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI909/MM11 N_WBLB<15>_XI909/MM11_d N_WWLB<7>_XI909/MM11_g
+ N_XI909/QB_XI909/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI909/MM1 N_XI909/Q_XI909/MM1_d N_XI909/QB_XI909/MM1_g N_GND_XI909/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI909/MM0 N_XI909/QB_XI909/MM0_d N_XI909/Q_XI909/MM0_g N_GND_XI909/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI909/MM9 N_XI909/NET08_XI909/MM9_d N_RWLB<7>_XI909/MM9_g N_RBL<15>_XI909/MM9_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI909/MM6 N_XI909/NET08_XI909/MM6_d N_XI909/QB_XI909/MM6_g N_VDD_XI909/MM6_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI909/MM5 N_XI909/Q_XI909/MM5_d N_XI909/QB_XI909/MM5_g N_VDD_XI909/MM5_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI909/MM4 N_XI909/QB_XI909/MM4_d N_XI909/Q_XI909/MM4_g N_VDD_XI909/MM4_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI908/MM8 N_XI908/NET08_XI908/MM8_d N_RWL<7>_XI908/MM8_g N_RBL<0>_XI908/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI908/MM7 N_XI908/NET08_XI908/MM7_d N_XI908/QB_XI908/MM7_g N_GND_XI908/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI908/MM10 N_WBL<0>_XI908/MM10_d N_WWLB<7>_XI908/MM10_g N_XI908/Q_XI908/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI908/MM11 N_WBLB<0>_XI908/MM11_d N_WWLB<7>_XI908/MM11_g
+ N_XI908/QB_XI908/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI908/MM1 N_XI908/Q_XI908/MM1_d N_XI908/QB_XI908/MM1_g N_GND_XI908/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI908/MM0 N_XI908/QB_XI908/MM0_d N_XI908/Q_XI908/MM0_g N_GND_XI908/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI908/MM9 N_XI908/NET08_XI908/MM9_d N_RWLB<7>_XI908/MM9_g N_RBL<0>_XI908/MM9_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI908/MM6 N_XI908/NET08_XI908/MM6_d N_XI908/QB_XI908/MM6_g N_VDD_XI908/MM6_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI908/MM5 N_XI908/Q_XI908/MM5_d N_XI908/QB_XI908/MM5_g N_VDD_XI908/MM5_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI908/MM4 N_XI908/QB_XI908/MM4_d N_XI908/Q_XI908/MM4_g N_VDD_XI908/MM4_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI907/MM8 N_XI907/NET08_XI907/MM8_d N_RWL<7>_XI907/MM8_g N_RBL<1>_XI907/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI907/MM7 N_XI907/NET08_XI907/MM7_d N_XI907/QB_XI907/MM7_g N_GND_XI907/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI907/MM10 N_WBL<1>_XI907/MM10_d N_WWLB<7>_XI907/MM10_g N_XI907/Q_XI907/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI907/MM11 N_WBLB<1>_XI907/MM11_d N_WWLB<7>_XI907/MM11_g
+ N_XI907/QB_XI907/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI907/MM1 N_XI907/Q_XI907/MM1_d N_XI907/QB_XI907/MM1_g N_GND_XI907/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI907/MM0 N_XI907/QB_XI907/MM0_d N_XI907/Q_XI907/MM0_g N_GND_XI907/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI907/MM9 N_XI907/NET08_XI907/MM9_d N_RWLB<7>_XI907/MM9_g N_RBL<1>_XI907/MM9_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI907/MM6 N_XI907/NET08_XI907/MM6_d N_XI907/QB_XI907/MM6_g N_VDD_XI907/MM6_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI907/MM5 N_XI907/Q_XI907/MM5_d N_XI907/QB_XI907/MM5_g N_VDD_XI907/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI907/MM4 N_XI907/QB_XI907/MM4_d N_XI907/Q_XI907/MM4_g N_VDD_XI907/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI906/MM8 N_XI906/NET08_XI906/MM8_d N_RWL<7>_XI906/MM8_g N_RBL<2>_XI906/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI906/MM7 N_XI906/NET08_XI906/MM7_d N_XI906/QB_XI906/MM7_g N_GND_XI906/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI906/MM10 N_WBL<2>_XI906/MM10_d N_WWLB<7>_XI906/MM10_g N_XI906/Q_XI906/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI906/MM11 N_WBLB<2>_XI906/MM11_d N_WWLB<7>_XI906/MM11_g
+ N_XI906/QB_XI906/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI906/MM1 N_XI906/Q_XI906/MM1_d N_XI906/QB_XI906/MM1_g N_GND_XI906/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI906/MM0 N_XI906/QB_XI906/MM0_d N_XI906/Q_XI906/MM0_g N_GND_XI906/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI906/MM9 N_XI906/NET08_XI906/MM9_d N_RWLB<7>_XI906/MM9_g N_RBL<2>_XI906/MM9_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI906/MM6 N_XI906/NET08_XI906/MM6_d N_XI906/QB_XI906/MM6_g N_VDD_XI906/MM6_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI906/MM5 N_XI906/Q_XI906/MM5_d N_XI906/QB_XI906/MM5_g N_VDD_XI906/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI906/MM4 N_XI906/QB_XI906/MM4_d N_XI906/Q_XI906/MM4_g N_VDD_XI906/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI895/MM8 N_XI895/NET08_XI895/MM8_d N_RWL<7>_XI895/MM8_g N_RBL<13>_XI895/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI895/MM7 N_XI895/NET08_XI895/MM7_d N_XI895/QB_XI895/MM7_g N_GND_XI895/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI895/MM10 N_WBL<13>_XI895/MM10_d N_WWLB<7>_XI895/MM10_g N_XI895/Q_XI895/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI895/MM11 N_WBLB<13>_XI895/MM11_d N_WWLB<7>_XI895/MM11_g
+ N_XI895/QB_XI895/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI895/MM1 N_XI895/Q_XI895/MM1_d N_XI895/QB_XI895/MM1_g N_GND_XI895/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI895/MM0 N_XI895/QB_XI895/MM0_d N_XI895/Q_XI895/MM0_g N_GND_XI895/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI895/MM9 N_XI895/NET08_XI895/MM9_d N_RWLB<7>_XI895/MM9_g N_RBL<13>_XI895/MM9_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI895/MM6 N_XI895/NET08_XI895/MM6_d N_XI895/QB_XI895/MM6_g N_VDD_XI895/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI895/MM5 N_XI895/Q_XI895/MM5_d N_XI895/QB_XI895/MM5_g N_VDD_XI895/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI895/MM4 N_XI895/QB_XI895/MM4_d N_XI895/Q_XI895/MM4_g N_VDD_XI895/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI894/MM8 N_XI894/NET08_XI894/MM8_d N_RWL<7>_XI894/MM8_g N_RBL<14>_XI894/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI894/MM7 N_XI894/NET08_XI894/MM7_d N_XI894/QB_XI894/MM7_g N_GND_XI894/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI894/MM10 N_WBL<14>_XI894/MM10_d N_WWLB<7>_XI894/MM10_g N_XI894/Q_XI894/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI894/MM11 N_WBLB<14>_XI894/MM11_d N_WWLB<7>_XI894/MM11_g
+ N_XI894/QB_XI894/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI894/MM1 N_XI894/Q_XI894/MM1_d N_XI894/QB_XI894/MM1_g N_GND_XI894/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI894/MM0 N_XI894/QB_XI894/MM0_d N_XI894/Q_XI894/MM0_g N_GND_XI894/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI894/MM9 N_XI894/NET08_XI894/MM9_d N_RWLB<7>_XI894/MM9_g N_RBL<14>_XI894/MM9_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI894/MM6 N_XI894/NET08_XI894/MM6_d N_XI894/QB_XI894/MM6_g N_VDD_XI894/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI894/MM5 N_XI894/Q_XI894/MM5_d N_XI894/QB_XI894/MM5_g N_VDD_XI894/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI894/MM4 N_XI894/QB_XI894/MM4_d N_XI894/Q_XI894/MM4_g N_VDD_XI894/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI927/MM8 N_XI927/NET08_XI927/MM8_d N_RWL<9>_XI927/MM8_g N_RBL<13>_XI927/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI927/MM7 N_XI927/NET08_XI927/MM7_d N_XI927/QB_XI927/MM7_g N_GND_XI927/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI927/MM10 N_WBL<13>_XI927/MM10_d N_WWLB<9>_XI927/MM10_g N_XI927/Q_XI927/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI927/MM11 N_WBLB<13>_XI927/MM11_d N_WWLB<9>_XI927/MM11_g
+ N_XI927/QB_XI927/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI927/MM1 N_XI927/Q_XI927/MM1_d N_XI927/QB_XI927/MM1_g N_GND_XI927/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI927/MM0 N_XI927/QB_XI927/MM0_d N_XI927/Q_XI927/MM0_g N_GND_XI927/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI927/MM9 N_XI927/NET08_XI927/MM9_d N_RWLB<9>_XI927/MM9_g N_RBL<13>_XI927/MM9_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI927/MM6 N_XI927/NET08_XI927/MM6_d N_XI927/QB_XI927/MM6_g N_VDD_XI927/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI927/MM5 N_XI927/Q_XI927/MM5_d N_XI927/QB_XI927/MM5_g N_VDD_XI927/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI927/MM4 N_XI927/QB_XI927/MM4_d N_XI927/Q_XI927/MM4_g N_VDD_XI927/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI926/MM8 N_XI926/NET08_XI926/MM8_d N_RWL<9>_XI926/MM8_g N_RBL<14>_XI926/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI926/MM7 N_XI926/NET08_XI926/MM7_d N_XI926/QB_XI926/MM7_g N_GND_XI926/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI926/MM10 N_WBL<14>_XI926/MM10_d N_WWLB<9>_XI926/MM10_g N_XI926/Q_XI926/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI926/MM11 N_WBLB<14>_XI926/MM11_d N_WWLB<9>_XI926/MM11_g
+ N_XI926/QB_XI926/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI926/MM1 N_XI926/Q_XI926/MM1_d N_XI926/QB_XI926/MM1_g N_GND_XI926/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI926/MM0 N_XI926/QB_XI926/MM0_d N_XI926/Q_XI926/MM0_g N_GND_XI926/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI926/MM9 N_XI926/NET08_XI926/MM9_d N_RWLB<9>_XI926/MM9_g N_RBL<14>_XI926/MM9_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI926/MM6 N_XI926/NET08_XI926/MM6_d N_XI926/QB_XI926/MM6_g N_VDD_XI926/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI926/MM5 N_XI926/Q_XI926/MM5_d N_XI926/QB_XI926/MM5_g N_VDD_XI926/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI926/MM4 N_XI926/QB_XI926/MM4_d N_XI926/Q_XI926/MM4_g N_VDD_XI926/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI925/MM8 N_XI925/NET08_XI925/MM8_d N_RWL<8>_XI925/MM8_g N_RBL<15>_XI925/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI925/MM7 N_XI925/NET08_XI925/MM7_d N_XI925/QB_XI925/MM7_g N_GND_XI925/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI925/MM10 N_WBL<15>_XI925/MM10_d N_WWLB<8>_XI925/MM10_g N_XI925/Q_XI925/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI925/MM11 N_WBLB<15>_XI925/MM11_d N_WWLB<8>_XI925/MM11_g
+ N_XI925/QB_XI925/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI925/MM1 N_XI925/Q_XI925/MM1_d N_XI925/QB_XI925/MM1_g N_GND_XI925/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI925/MM0 N_XI925/QB_XI925/MM0_d N_XI925/Q_XI925/MM0_g N_GND_XI925/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI925/MM9 N_XI925/NET08_XI925/MM9_d N_RWLB<8>_XI925/MM9_g N_RBL<15>_XI925/MM9_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI925/MM6 N_XI925/NET08_XI925/MM6_d N_XI925/QB_XI925/MM6_g N_VDD_XI925/MM6_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI925/MM5 N_XI925/Q_XI925/MM5_d N_XI925/QB_XI925/MM5_g N_VDD_XI925/MM5_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI925/MM4 N_XI925/QB_XI925/MM4_d N_XI925/Q_XI925/MM4_g N_VDD_XI925/MM4_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI924/MM8 N_XI924/NET08_XI924/MM8_d N_RWL<8>_XI924/MM8_g N_RBL<0>_XI924/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI924/MM7 N_XI924/NET08_XI924/MM7_d N_XI924/QB_XI924/MM7_g N_GND_XI924/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI924/MM10 N_WBL<0>_XI924/MM10_d N_WWLB<8>_XI924/MM10_g N_XI924/Q_XI924/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI924/MM11 N_WBLB<0>_XI924/MM11_d N_WWLB<8>_XI924/MM11_g
+ N_XI924/QB_XI924/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI924/MM1 N_XI924/Q_XI924/MM1_d N_XI924/QB_XI924/MM1_g N_GND_XI924/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI924/MM0 N_XI924/QB_XI924/MM0_d N_XI924/Q_XI924/MM0_g N_GND_XI924/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI924/MM9 N_XI924/NET08_XI924/MM9_d N_RWLB<8>_XI924/MM9_g N_RBL<0>_XI924/MM9_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI924/MM6 N_XI924/NET08_XI924/MM6_d N_XI924/QB_XI924/MM6_g N_VDD_XI924/MM6_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI924/MM5 N_XI924/Q_XI924/MM5_d N_XI924/QB_XI924/MM5_g N_VDD_XI924/MM5_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI924/MM4 N_XI924/QB_XI924/MM4_d N_XI924/Q_XI924/MM4_g N_VDD_XI924/MM4_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1030/MM8 N_XI1030/NET08_XI1030/MM8_d N_RWL<15>_XI1030/MM8_g
+ N_RBL<6>_XI1030/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1030/MM7 N_XI1030/NET08_XI1030/MM7_d N_XI1030/QB_XI1030/MM7_g
+ N_GND_XI1030/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1030/MM10 N_WBL<6>_XI1030/MM10_d N_WWLB<15>_XI1030/MM10_g
+ N_XI1030/Q_XI1030/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1030/MM11 N_WBLB<6>_XI1030/MM11_d N_WWLB<15>_XI1030/MM11_g
+ N_XI1030/QB_XI1030/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1030/MM1 N_XI1030/Q_XI1030/MM1_d N_XI1030/QB_XI1030/MM1_g N_GND_XI1030/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1030/MM0 N_XI1030/QB_XI1030/MM0_d N_XI1030/Q_XI1030/MM0_g N_GND_XI1030/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1030/MM9 N_XI1030/NET08_XI1030/MM9_d N_RWLB<15>_XI1030/MM9_g
+ N_RBL<6>_XI1030/MM9_s N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1030/MM6 N_XI1030/NET08_XI1030/MM6_d N_XI1030/QB_XI1030/MM6_g
+ N_VDD_XI1030/MM6_s N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1030/MM5 N_XI1030/Q_XI1030/MM5_d N_XI1030/QB_XI1030/MM5_g N_VDD_XI1030/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1030/MM4 N_XI1030/QB_XI1030/MM4_d N_XI1030/Q_XI1030/MM4_g N_VDD_XI1030/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI997/MM8 N_XI997/NET08_XI997/MM8_d N_RWL<13>_XI997/MM8_g N_RBL<7>_XI997/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI997/MM7 N_XI997/NET08_XI997/MM7_d N_XI997/QB_XI997/MM7_g N_GND_XI997/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI997/MM10 N_WBL<7>_XI997/MM10_d N_WWLB<13>_XI997/MM10_g N_XI997/Q_XI997/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI997/MM11 N_WBLB<7>_XI997/MM11_d N_WWLB<13>_XI997/MM11_g
+ N_XI997/QB_XI997/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI997/MM1 N_XI997/Q_XI997/MM1_d N_XI997/QB_XI997/MM1_g N_GND_XI997/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI997/MM0 N_XI997/QB_XI997/MM0_d N_XI997/Q_XI997/MM0_g N_GND_XI997/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI997/MM9 N_XI997/NET08_XI997/MM9_d N_RWLB<13>_XI997/MM9_g N_RBL<7>_XI997/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI997/MM6 N_XI997/NET08_XI997/MM6_d N_XI997/QB_XI997/MM6_g N_VDD_XI997/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI997/MM5 N_XI997/Q_XI997/MM5_d N_XI997/QB_XI997/MM5_g N_VDD_XI997/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI997/MM4 N_XI997/QB_XI997/MM4_d N_XI997/Q_XI997/MM4_g N_VDD_XI997/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI871/MM8 N_XI871/NET08_XI871/MM8_d N_RWL<5>_XI871/MM8_g N_RBL<5>_XI871/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI871/MM7 N_XI871/NET08_XI871/MM7_d N_XI871/QB_XI871/MM7_g N_GND_XI871/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI871/MM10 N_WBL<5>_XI871/MM10_d N_WWLB<5>_XI871/MM10_g N_XI871/Q_XI871/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI871/MM11 N_WBLB<5>_XI871/MM11_d N_WWLB<5>_XI871/MM11_g
+ N_XI871/QB_XI871/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI871/MM1 N_XI871/Q_XI871/MM1_d N_XI871/QB_XI871/MM1_g N_GND_XI871/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI871/MM0 N_XI871/QB_XI871/MM0_d N_XI871/Q_XI871/MM0_g N_GND_XI871/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI871/MM9 N_XI871/NET08_XI871/MM9_d N_RWLB<5>_XI871/MM9_g N_RBL<5>_XI871/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI871/MM6 N_XI871/NET08_XI871/MM6_d N_XI871/QB_XI871/MM6_g N_VDD_XI871/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI871/MM5 N_XI871/Q_XI871/MM5_d N_XI871/QB_XI871/MM5_g N_VDD_XI871/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI871/MM4 N_XI871/QB_XI871/MM4_d N_XI871/Q_XI871/MM4_g N_VDD_XI871/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI870/MM8 N_XI870/NET08_XI870/MM8_d N_RWL<5>_XI870/MM8_g N_RBL<6>_XI870/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI870/MM7 N_XI870/NET08_XI870/MM7_d N_XI870/QB_XI870/MM7_g N_GND_XI870/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI870/MM10 N_WBL<6>_XI870/MM10_d N_WWLB<5>_XI870/MM10_g N_XI870/Q_XI870/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI870/MM11 N_WBLB<6>_XI870/MM11_d N_WWLB<5>_XI870/MM11_g
+ N_XI870/QB_XI870/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI870/MM1 N_XI870/Q_XI870/MM1_d N_XI870/QB_XI870/MM1_g N_GND_XI870/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI870/MM0 N_XI870/QB_XI870/MM0_d N_XI870/Q_XI870/MM0_g N_GND_XI870/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI870/MM9 N_XI870/NET08_XI870/MM9_d N_RWLB<5>_XI870/MM9_g N_RBL<6>_XI870/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI870/MM6 N_XI870/NET08_XI870/MM6_d N_XI870/QB_XI870/MM6_g N_VDD_XI870/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI870/MM5 N_XI870/Q_XI870/MM5_d N_XI870/QB_XI870/MM5_g N_VDD_XI870/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI870/MM4 N_XI870/QB_XI870/MM4_d N_XI870/Q_XI870/MM4_g N_VDD_XI870/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI869/MM8 N_XI869/NET08_XI869/MM8_d N_RWL<5>_XI869/MM8_g N_RBL<7>_XI869/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI869/MM7 N_XI869/NET08_XI869/MM7_d N_XI869/QB_XI869/MM7_g N_GND_XI869/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI869/MM10 N_WBL<7>_XI869/MM10_d N_WWLB<5>_XI869/MM10_g N_XI869/Q_XI869/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI869/MM11 N_WBLB<7>_XI869/MM11_d N_WWLB<5>_XI869/MM11_g
+ N_XI869/QB_XI869/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI869/MM1 N_XI869/Q_XI869/MM1_d N_XI869/QB_XI869/MM1_g N_GND_XI869/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI869/MM0 N_XI869/QB_XI869/MM0_d N_XI869/Q_XI869/MM0_g N_GND_XI869/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI869/MM9 N_XI869/NET08_XI869/MM9_d N_RWLB<5>_XI869/MM9_g N_RBL<7>_XI869/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI869/MM6 N_XI869/NET08_XI869/MM6_d N_XI869/QB_XI869/MM6_g N_VDD_XI869/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI869/MM5 N_XI869/Q_XI869/MM5_d N_XI869/QB_XI869/MM5_g N_VDD_XI869/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI869/MM4 N_XI869/QB_XI869/MM4_d N_XI869/Q_XI869/MM4_g N_VDD_XI869/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI868/MM8 N_XI868/NET08_XI868/MM8_d N_RWL<5>_XI868/MM8_g N_RBL<8>_XI868/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI868/MM7 N_XI868/NET08_XI868/MM7_d N_XI868/QB_XI868/MM7_g N_GND_XI868/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI868/MM10 N_WBL<8>_XI868/MM10_d N_WWLB<5>_XI868/MM10_g N_XI868/Q_XI868/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI868/MM11 N_WBLB<8>_XI868/MM11_d N_WWLB<5>_XI868/MM11_g
+ N_XI868/QB_XI868/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI868/MM1 N_XI868/Q_XI868/MM1_d N_XI868/QB_XI868/MM1_g N_GND_XI868/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI868/MM0 N_XI868/QB_XI868/MM0_d N_XI868/Q_XI868/MM0_g N_GND_XI868/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI868/MM9 N_XI868/NET08_XI868/MM9_d N_RWLB<5>_XI868/MM9_g N_RBL<8>_XI868/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI868/MM6 N_XI868/NET08_XI868/MM6_d N_XI868/QB_XI868/MM6_g N_VDD_XI868/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI868/MM5 N_XI868/Q_XI868/MM5_d N_XI868/QB_XI868/MM5_g N_VDD_XI868/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI868/MM4 N_XI868/QB_XI868/MM4_d N_XI868/Q_XI868/MM4_g N_VDD_XI868/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI905/MM8 N_XI905/NET08_XI905/MM8_d N_RWL<7>_XI905/MM8_g N_RBL<3>_XI905/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI905/MM7 N_XI905/NET08_XI905/MM7_d N_XI905/QB_XI905/MM7_g N_GND_XI905/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI905/MM10 N_WBL<3>_XI905/MM10_d N_WWLB<7>_XI905/MM10_g N_XI905/Q_XI905/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI905/MM11 N_WBLB<3>_XI905/MM11_d N_WWLB<7>_XI905/MM11_g
+ N_XI905/QB_XI905/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI905/MM1 N_XI905/Q_XI905/MM1_d N_XI905/QB_XI905/MM1_g N_GND_XI905/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI905/MM0 N_XI905/QB_XI905/MM0_d N_XI905/Q_XI905/MM0_g N_GND_XI905/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI905/MM9 N_XI905/NET08_XI905/MM9_d N_RWLB<7>_XI905/MM9_g N_RBL<3>_XI905/MM9_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI905/MM6 N_XI905/NET08_XI905/MM6_d N_XI905/QB_XI905/MM6_g N_VDD_XI905/MM6_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI905/MM5 N_XI905/Q_XI905/MM5_d N_XI905/QB_XI905/MM5_g N_VDD_XI905/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI905/MM4 N_XI905/QB_XI905/MM4_d N_XI905/Q_XI905/MM4_g N_VDD_XI905/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI904/MM8 N_XI904/NET08_XI904/MM8_d N_RWL<7>_XI904/MM8_g N_RBL<4>_XI904/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI904/MM7 N_XI904/NET08_XI904/MM7_d N_XI904/QB_XI904/MM7_g N_GND_XI904/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI904/MM10 N_WBL<4>_XI904/MM10_d N_WWLB<7>_XI904/MM10_g N_XI904/Q_XI904/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI904/MM11 N_WBLB<4>_XI904/MM11_d N_WWLB<7>_XI904/MM11_g
+ N_XI904/QB_XI904/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI904/MM1 N_XI904/Q_XI904/MM1_d N_XI904/QB_XI904/MM1_g N_GND_XI904/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI904/MM0 N_XI904/QB_XI904/MM0_d N_XI904/Q_XI904/MM0_g N_GND_XI904/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI904/MM9 N_XI904/NET08_XI904/MM9_d N_RWLB<7>_XI904/MM9_g N_RBL<4>_XI904/MM9_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI904/MM6 N_XI904/NET08_XI904/MM6_d N_XI904/QB_XI904/MM6_g N_VDD_XI904/MM6_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI904/MM5 N_XI904/Q_XI904/MM5_d N_XI904/QB_XI904/MM5_g N_VDD_XI904/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI904/MM4 N_XI904/QB_XI904/MM4_d N_XI904/Q_XI904/MM4_g N_VDD_XI904/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI903/MM8 N_XI903/NET08_XI903/MM8_d N_RWL<7>_XI903/MM8_g N_RBL<5>_XI903/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI903/MM7 N_XI903/NET08_XI903/MM7_d N_XI903/QB_XI903/MM7_g N_GND_XI903/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI903/MM10 N_WBL<5>_XI903/MM10_d N_WWLB<7>_XI903/MM10_g N_XI903/Q_XI903/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI903/MM11 N_WBLB<5>_XI903/MM11_d N_WWLB<7>_XI903/MM11_g
+ N_XI903/QB_XI903/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI903/MM1 N_XI903/Q_XI903/MM1_d N_XI903/QB_XI903/MM1_g N_GND_XI903/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI903/MM0 N_XI903/QB_XI903/MM0_d N_XI903/Q_XI903/MM0_g N_GND_XI903/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI903/MM9 N_XI903/NET08_XI903/MM9_d N_RWLB<7>_XI903/MM9_g N_RBL<5>_XI903/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI903/MM6 N_XI903/NET08_XI903/MM6_d N_XI903/QB_XI903/MM6_g N_VDD_XI903/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI903/MM5 N_XI903/Q_XI903/MM5_d N_XI903/QB_XI903/MM5_g N_VDD_XI903/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI903/MM4 N_XI903/QB_XI903/MM4_d N_XI903/Q_XI903/MM4_g N_VDD_XI903/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI902/MM8 N_XI902/NET08_XI902/MM8_d N_RWL<7>_XI902/MM8_g N_RBL<6>_XI902/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI902/MM7 N_XI902/NET08_XI902/MM7_d N_XI902/QB_XI902/MM7_g N_GND_XI902/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI902/MM10 N_WBL<6>_XI902/MM10_d N_WWLB<7>_XI902/MM10_g N_XI902/Q_XI902/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI902/MM11 N_WBLB<6>_XI902/MM11_d N_WWLB<7>_XI902/MM11_g
+ N_XI902/QB_XI902/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI902/MM1 N_XI902/Q_XI902/MM1_d N_XI902/QB_XI902/MM1_g N_GND_XI902/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI902/MM0 N_XI902/QB_XI902/MM0_d N_XI902/Q_XI902/MM0_g N_GND_XI902/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI902/MM9 N_XI902/NET08_XI902/MM9_d N_RWLB<7>_XI902/MM9_g N_RBL<6>_XI902/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI902/MM6 N_XI902/NET08_XI902/MM6_d N_XI902/QB_XI902/MM6_g N_VDD_XI902/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI902/MM5 N_XI902/Q_XI902/MM5_d N_XI902/QB_XI902/MM5_g N_VDD_XI902/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI902/MM4 N_XI902/QB_XI902/MM4_d N_XI902/Q_XI902/MM4_g N_VDD_XI902/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI901/MM8 N_XI901/NET08_XI901/MM8_d N_RWL<7>_XI901/MM8_g N_RBL<7>_XI901/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI901/MM7 N_XI901/NET08_XI901/MM7_d N_XI901/QB_XI901/MM7_g N_GND_XI901/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI901/MM10 N_WBL<7>_XI901/MM10_d N_WWLB<7>_XI901/MM10_g N_XI901/Q_XI901/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI901/MM11 N_WBLB<7>_XI901/MM11_d N_WWLB<7>_XI901/MM11_g
+ N_XI901/QB_XI901/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI901/MM1 N_XI901/Q_XI901/MM1_d N_XI901/QB_XI901/MM1_g N_GND_XI901/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI901/MM0 N_XI901/QB_XI901/MM0_d N_XI901/Q_XI901/MM0_g N_GND_XI901/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI901/MM9 N_XI901/NET08_XI901/MM9_d N_RWLB<7>_XI901/MM9_g N_RBL<7>_XI901/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI901/MM6 N_XI901/NET08_XI901/MM6_d N_XI901/QB_XI901/MM6_g N_VDD_XI901/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI901/MM5 N_XI901/Q_XI901/MM5_d N_XI901/QB_XI901/MM5_g N_VDD_XI901/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI901/MM4 N_XI901/QB_XI901/MM4_d N_XI901/Q_XI901/MM4_g N_VDD_XI901/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI890/MM8 N_XI890/NET08_XI890/MM8_d N_RWL<6>_XI890/MM8_g N_RBL<2>_XI890/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI890/MM7 N_XI890/NET08_XI890/MM7_d N_XI890/QB_XI890/MM7_g N_GND_XI890/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI890/MM10 N_WBL<2>_XI890/MM10_d N_WWLB<6>_XI890/MM10_g N_XI890/Q_XI890/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI890/MM11 N_WBLB<2>_XI890/MM11_d N_WWLB<6>_XI890/MM11_g
+ N_XI890/QB_XI890/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI890/MM1 N_XI890/Q_XI890/MM1_d N_XI890/QB_XI890/MM1_g N_GND_XI890/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI890/MM0 N_XI890/QB_XI890/MM0_d N_XI890/Q_XI890/MM0_g N_GND_XI890/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI890/MM9 N_XI890/NET08_XI890/MM9_d N_RWLB<6>_XI890/MM9_g N_RBL<2>_XI890/MM9_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI890/MM6 N_XI890/NET08_XI890/MM6_d N_XI890/QB_XI890/MM6_g N_VDD_XI890/MM6_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI890/MM5 N_XI890/Q_XI890/MM5_d N_XI890/QB_XI890/MM5_g N_VDD_XI890/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI890/MM4 N_XI890/QB_XI890/MM4_d N_XI890/Q_XI890/MM4_g N_VDD_XI890/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI889/MM8 N_XI889/NET08_XI889/MM8_d N_RWL<6>_XI889/MM8_g N_RBL<3>_XI889/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI889/MM7 N_XI889/NET08_XI889/MM7_d N_XI889/QB_XI889/MM7_g N_GND_XI889/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI889/MM10 N_WBL<3>_XI889/MM10_d N_WWLB<6>_XI889/MM10_g N_XI889/Q_XI889/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI889/MM11 N_WBLB<3>_XI889/MM11_d N_WWLB<6>_XI889/MM11_g
+ N_XI889/QB_XI889/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI889/MM1 N_XI889/Q_XI889/MM1_d N_XI889/QB_XI889/MM1_g N_GND_XI889/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI889/MM0 N_XI889/QB_XI889/MM0_d N_XI889/Q_XI889/MM0_g N_GND_XI889/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI889/MM9 N_XI889/NET08_XI889/MM9_d N_RWLB<6>_XI889/MM9_g N_RBL<3>_XI889/MM9_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI889/MM6 N_XI889/NET08_XI889/MM6_d N_XI889/QB_XI889/MM6_g N_VDD_XI889/MM6_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI889/MM5 N_XI889/Q_XI889/MM5_d N_XI889/QB_XI889/MM5_g N_VDD_XI889/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI889/MM4 N_XI889/QB_XI889/MM4_d N_XI889/Q_XI889/MM4_g N_VDD_XI889/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI888/MM8 N_XI888/NET08_XI888/MM8_d N_RWL<6>_XI888/MM8_g N_RBL<4>_XI888/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI888/MM7 N_XI888/NET08_XI888/MM7_d N_XI888/QB_XI888/MM7_g N_GND_XI888/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI888/MM10 N_WBL<4>_XI888/MM10_d N_WWLB<6>_XI888/MM10_g N_XI888/Q_XI888/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI888/MM11 N_WBLB<4>_XI888/MM11_d N_WWLB<6>_XI888/MM11_g
+ N_XI888/QB_XI888/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI888/MM1 N_XI888/Q_XI888/MM1_d N_XI888/QB_XI888/MM1_g N_GND_XI888/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI888/MM0 N_XI888/QB_XI888/MM0_d N_XI888/Q_XI888/MM0_g N_GND_XI888/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI888/MM9 N_XI888/NET08_XI888/MM9_d N_RWLB<6>_XI888/MM9_g N_RBL<4>_XI888/MM9_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI888/MM6 N_XI888/NET08_XI888/MM6_d N_XI888/QB_XI888/MM6_g N_VDD_XI888/MM6_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI888/MM5 N_XI888/Q_XI888/MM5_d N_XI888/QB_XI888/MM5_g N_VDD_XI888/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI888/MM4 N_XI888/QB_XI888/MM4_d N_XI888/Q_XI888/MM4_g N_VDD_XI888/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI923/MM8 N_XI923/NET08_XI923/MM8_d N_RWL<8>_XI923/MM8_g N_RBL<1>_XI923/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI923/MM7 N_XI923/NET08_XI923/MM7_d N_XI923/QB_XI923/MM7_g N_GND_XI923/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI923/MM10 N_WBL<1>_XI923/MM10_d N_WWLB<8>_XI923/MM10_g N_XI923/Q_XI923/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI923/MM11 N_WBLB<1>_XI923/MM11_d N_WWLB<8>_XI923/MM11_g
+ N_XI923/QB_XI923/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI923/MM1 N_XI923/Q_XI923/MM1_d N_XI923/QB_XI923/MM1_g N_GND_XI923/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI923/MM0 N_XI923/QB_XI923/MM0_d N_XI923/Q_XI923/MM0_g N_GND_XI923/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI923/MM9 N_XI923/NET08_XI923/MM9_d N_RWLB<8>_XI923/MM9_g N_RBL<1>_XI923/MM9_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI923/MM6 N_XI923/NET08_XI923/MM6_d N_XI923/QB_XI923/MM6_g N_VDD_XI923/MM6_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI923/MM5 N_XI923/Q_XI923/MM5_d N_XI923/QB_XI923/MM5_g N_VDD_XI923/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI923/MM4 N_XI923/QB_XI923/MM4_d N_XI923/Q_XI923/MM4_g N_VDD_XI923/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI922/MM8 N_XI922/NET08_XI922/MM8_d N_RWL<8>_XI922/MM8_g N_RBL<2>_XI922/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI922/MM7 N_XI922/NET08_XI922/MM7_d N_XI922/QB_XI922/MM7_g N_GND_XI922/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI922/MM10 N_WBL<2>_XI922/MM10_d N_WWLB<8>_XI922/MM10_g N_XI922/Q_XI922/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI922/MM11 N_WBLB<2>_XI922/MM11_d N_WWLB<8>_XI922/MM11_g
+ N_XI922/QB_XI922/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI922/MM1 N_XI922/Q_XI922/MM1_d N_XI922/QB_XI922/MM1_g N_GND_XI922/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI922/MM0 N_XI922/QB_XI922/MM0_d N_XI922/Q_XI922/MM0_g N_GND_XI922/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI922/MM9 N_XI922/NET08_XI922/MM9_d N_RWLB<8>_XI922/MM9_g N_RBL<2>_XI922/MM9_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI922/MM6 N_XI922/NET08_XI922/MM6_d N_XI922/QB_XI922/MM6_g N_VDD_XI922/MM6_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI922/MM5 N_XI922/Q_XI922/MM5_d N_XI922/QB_XI922/MM5_g N_VDD_XI922/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI922/MM4 N_XI922/QB_XI922/MM4_d N_XI922/Q_XI922/MM4_g N_VDD_XI922/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI921/MM8 N_XI921/NET08_XI921/MM8_d N_RWL<8>_XI921/MM8_g N_RBL<3>_XI921/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI921/MM7 N_XI921/NET08_XI921/MM7_d N_XI921/QB_XI921/MM7_g N_GND_XI921/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI921/MM10 N_WBL<3>_XI921/MM10_d N_WWLB<8>_XI921/MM10_g N_XI921/Q_XI921/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI921/MM11 N_WBLB<3>_XI921/MM11_d N_WWLB<8>_XI921/MM11_g
+ N_XI921/QB_XI921/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI921/MM1 N_XI921/Q_XI921/MM1_d N_XI921/QB_XI921/MM1_g N_GND_XI921/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI921/MM0 N_XI921/QB_XI921/MM0_d N_XI921/Q_XI921/MM0_g N_GND_XI921/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI921/MM9 N_XI921/NET08_XI921/MM9_d N_RWLB<8>_XI921/MM9_g N_RBL<3>_XI921/MM9_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI921/MM6 N_XI921/NET08_XI921/MM6_d N_XI921/QB_XI921/MM6_g N_VDD_XI921/MM6_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI921/MM5 N_XI921/Q_XI921/MM5_d N_XI921/QB_XI921/MM5_g N_VDD_XI921/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI921/MM4 N_XI921/QB_XI921/MM4_d N_XI921/Q_XI921/MM4_g N_VDD_XI921/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI920/MM8 N_XI920/NET08_XI920/MM8_d N_RWL<8>_XI920/MM8_g N_RBL<4>_XI920/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI920/MM7 N_XI920/NET08_XI920/MM7_d N_XI920/QB_XI920/MM7_g N_GND_XI920/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI920/MM10 N_WBL<4>_XI920/MM10_d N_WWLB<8>_XI920/MM10_g N_XI920/Q_XI920/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI920/MM11 N_WBLB<4>_XI920/MM11_d N_WWLB<8>_XI920/MM11_g
+ N_XI920/QB_XI920/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI920/MM1 N_XI920/Q_XI920/MM1_d N_XI920/QB_XI920/MM1_g N_GND_XI920/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI920/MM0 N_XI920/QB_XI920/MM0_d N_XI920/Q_XI920/MM0_g N_GND_XI920/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI920/MM9 N_XI920/NET08_XI920/MM9_d N_RWLB<8>_XI920/MM9_g N_RBL<4>_XI920/MM9_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI920/MM6 N_XI920/NET08_XI920/MM6_d N_XI920/QB_XI920/MM6_g N_VDD_XI920/MM6_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI920/MM5 N_XI920/Q_XI920/MM5_d N_XI920/QB_XI920/MM5_g N_VDD_XI920/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI920/MM4 N_XI920/QB_XI920/MM4_d N_XI920/Q_XI920/MM4_g N_VDD_XI920/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1029/MM8 N_XI1029/NET08_XI1029/MM8_d N_RWL<15>_XI1029/MM8_g
+ N_RBL<7>_XI1029/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1029/MM7 N_XI1029/NET08_XI1029/MM7_d N_XI1029/QB_XI1029/MM7_g
+ N_GND_XI1029/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1029/MM10 N_WBL<7>_XI1029/MM10_d N_WWLB<15>_XI1029/MM10_g
+ N_XI1029/Q_XI1029/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1029/MM11 N_WBLB<7>_XI1029/MM11_d N_WWLB<15>_XI1029/MM11_g
+ N_XI1029/QB_XI1029/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1029/MM1 N_XI1029/Q_XI1029/MM1_d N_XI1029/QB_XI1029/MM1_g N_GND_XI1029/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1029/MM0 N_XI1029/QB_XI1029/MM0_d N_XI1029/Q_XI1029/MM0_g N_GND_XI1029/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1029/MM9 N_XI1029/NET08_XI1029/MM9_d N_RWLB<15>_XI1029/MM9_g
+ N_RBL<7>_XI1029/MM9_s N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1029/MM6 N_XI1029/NET08_XI1029/MM6_d N_XI1029/QB_XI1029/MM6_g
+ N_VDD_XI1029/MM6_s N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1029/MM5 N_XI1029/Q_XI1029/MM5_d N_XI1029/QB_XI1029/MM5_g N_VDD_XI1029/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1029/MM4 N_XI1029/QB_XI1029/MM4_d N_XI1029/Q_XI1029/MM4_g N_VDD_XI1029/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI998/MM8 N_XI998/NET08_XI998/MM8_d N_RWL<13>_XI998/MM8_g N_RBL<6>_XI998/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI998/MM7 N_XI998/NET08_XI998/MM7_d N_XI998/QB_XI998/MM7_g N_GND_XI998/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI998/MM10 N_WBL<6>_XI998/MM10_d N_WWLB<13>_XI998/MM10_g N_XI998/Q_XI998/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI998/MM11 N_WBLB<6>_XI998/MM11_d N_WWLB<13>_XI998/MM11_g
+ N_XI998/QB_XI998/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI998/MM1 N_XI998/Q_XI998/MM1_d N_XI998/QB_XI998/MM1_g N_GND_XI998/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI998/MM0 N_XI998/QB_XI998/MM0_d N_XI998/Q_XI998/MM0_g N_GND_XI998/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI998/MM9 N_XI998/NET08_XI998/MM9_d N_RWLB<13>_XI998/MM9_g N_RBL<6>_XI998/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI998/MM6 N_XI998/NET08_XI998/MM6_d N_XI998/QB_XI998/MM6_g N_VDD_XI998/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI998/MM5 N_XI998/Q_XI998/MM5_d N_XI998/QB_XI998/MM5_g N_VDD_XI998/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI998/MM4 N_XI998/QB_XI998/MM4_d N_XI998/Q_XI998/MM4_g N_VDD_XI998/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI867/MM8 N_XI867/NET08_XI867/MM8_d N_RWL<5>_XI867/MM8_g N_RBL<9>_XI867/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI867/MM7 N_XI867/NET08_XI867/MM7_d N_XI867/QB_XI867/MM7_g N_GND_XI867/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI867/MM10 N_WBL<9>_XI867/MM10_d N_WWLB<5>_XI867/MM10_g N_XI867/Q_XI867/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI867/MM11 N_WBLB<9>_XI867/MM11_d N_WWLB<5>_XI867/MM11_g
+ N_XI867/QB_XI867/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI867/MM1 N_XI867/Q_XI867/MM1_d N_XI867/QB_XI867/MM1_g N_GND_XI867/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI867/MM0 N_XI867/QB_XI867/MM0_d N_XI867/Q_XI867/MM0_g N_GND_XI867/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI867/MM9 N_XI867/NET08_XI867/MM9_d N_RWLB<5>_XI867/MM9_g N_RBL<9>_XI867/MM9_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI867/MM6 N_XI867/NET08_XI867/MM6_d N_XI867/QB_XI867/MM6_g N_VDD_XI867/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI867/MM5 N_XI867/Q_XI867/MM5_d N_XI867/QB_XI867/MM5_g N_VDD_XI867/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI867/MM4 N_XI867/QB_XI867/MM4_d N_XI867/Q_XI867/MM4_g N_VDD_XI867/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI866/MM8 N_XI866/NET08_XI866/MM8_d N_RWL<5>_XI866/MM8_g N_RBL<10>_XI866/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI866/MM7 N_XI866/NET08_XI866/MM7_d N_XI866/QB_XI866/MM7_g N_GND_XI866/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI866/MM10 N_WBL<10>_XI866/MM10_d N_WWLB<5>_XI866/MM10_g N_XI866/Q_XI866/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI866/MM11 N_WBLB<10>_XI866/MM11_d N_WWLB<5>_XI866/MM11_g
+ N_XI866/QB_XI866/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI866/MM1 N_XI866/Q_XI866/MM1_d N_XI866/QB_XI866/MM1_g N_GND_XI866/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI866/MM0 N_XI866/QB_XI866/MM0_d N_XI866/Q_XI866/MM0_g N_GND_XI866/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI866/MM9 N_XI866/NET08_XI866/MM9_d N_RWLB<5>_XI866/MM9_g N_RBL<10>_XI866/MM9_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI866/MM6 N_XI866/NET08_XI866/MM6_d N_XI866/QB_XI866/MM6_g N_VDD_XI866/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI866/MM5 N_XI866/Q_XI866/MM5_d N_XI866/QB_XI866/MM5_g N_VDD_XI866/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI866/MM4 N_XI866/QB_XI866/MM4_d N_XI866/Q_XI866/MM4_g N_VDD_XI866/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI865/MM8 N_XI865/NET08_XI865/MM8_d N_RWL<5>_XI865/MM8_g N_RBL<11>_XI865/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI865/MM7 N_XI865/NET08_XI865/MM7_d N_XI865/QB_XI865/MM7_g N_GND_XI865/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI865/MM10 N_WBL<11>_XI865/MM10_d N_WWLB<5>_XI865/MM10_g N_XI865/Q_XI865/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI865/MM11 N_WBLB<11>_XI865/MM11_d N_WWLB<5>_XI865/MM11_g
+ N_XI865/QB_XI865/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI865/MM1 N_XI865/Q_XI865/MM1_d N_XI865/QB_XI865/MM1_g N_GND_XI865/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI865/MM0 N_XI865/QB_XI865/MM0_d N_XI865/Q_XI865/MM0_g N_GND_XI865/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI865/MM9 N_XI865/NET08_XI865/MM9_d N_RWLB<5>_XI865/MM9_g N_RBL<11>_XI865/MM9_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI865/MM6 N_XI865/NET08_XI865/MM6_d N_XI865/QB_XI865/MM6_g N_VDD_XI865/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI865/MM5 N_XI865/Q_XI865/MM5_d N_XI865/QB_XI865/MM5_g N_VDD_XI865/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI865/MM4 N_XI865/QB_XI865/MM4_d N_XI865/Q_XI865/MM4_g N_VDD_XI865/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI864/MM8 N_XI864/NET08_XI864/MM8_d N_RWL<5>_XI864/MM8_g N_RBL<12>_XI864/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI864/MM7 N_XI864/NET08_XI864/MM7_d N_XI864/QB_XI864/MM7_g N_GND_XI864/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI864/MM10 N_WBL<12>_XI864/MM10_d N_WWLB<5>_XI864/MM10_g N_XI864/Q_XI864/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI864/MM11 N_WBLB<12>_XI864/MM11_d N_WWLB<5>_XI864/MM11_g
+ N_XI864/QB_XI864/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI864/MM1 N_XI864/Q_XI864/MM1_d N_XI864/QB_XI864/MM1_g N_GND_XI864/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI864/MM0 N_XI864/QB_XI864/MM0_d N_XI864/Q_XI864/MM0_g N_GND_XI864/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI864/MM9 N_XI864/NET08_XI864/MM9_d N_RWLB<5>_XI864/MM9_g N_RBL<12>_XI864/MM9_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI864/MM6 N_XI864/NET08_XI864/MM6_d N_XI864/QB_XI864/MM6_g N_VDD_XI864/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI864/MM5 N_XI864/Q_XI864/MM5_d N_XI864/QB_XI864/MM5_g N_VDD_XI864/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI864/MM4 N_XI864/QB_XI864/MM4_d N_XI864/Q_XI864/MM4_g N_VDD_XI864/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI899/MM8 N_XI899/NET08_XI899/MM8_d N_RWL<7>_XI899/MM8_g N_RBL<9>_XI899/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI899/MM7 N_XI899/NET08_XI899/MM7_d N_XI899/QB_XI899/MM7_g N_GND_XI899/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI899/MM10 N_WBL<9>_XI899/MM10_d N_WWLB<7>_XI899/MM10_g N_XI899/Q_XI899/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI899/MM11 N_WBLB<9>_XI899/MM11_d N_WWLB<7>_XI899/MM11_g
+ N_XI899/QB_XI899/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI899/MM1 N_XI899/Q_XI899/MM1_d N_XI899/QB_XI899/MM1_g N_GND_XI899/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI899/MM0 N_XI899/QB_XI899/MM0_d N_XI899/Q_XI899/MM0_g N_GND_XI899/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI899/MM9 N_XI899/NET08_XI899/MM9_d N_RWLB<7>_XI899/MM9_g N_RBL<9>_XI899/MM9_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI899/MM6 N_XI899/NET08_XI899/MM6_d N_XI899/QB_XI899/MM6_g N_VDD_XI899/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI899/MM5 N_XI899/Q_XI899/MM5_d N_XI899/QB_XI899/MM5_g N_VDD_XI899/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI899/MM4 N_XI899/QB_XI899/MM4_d N_XI899/Q_XI899/MM4_g N_VDD_XI899/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI898/MM8 N_XI898/NET08_XI898/MM8_d N_RWL<7>_XI898/MM8_g N_RBL<10>_XI898/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI898/MM7 N_XI898/NET08_XI898/MM7_d N_XI898/QB_XI898/MM7_g N_GND_XI898/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI898/MM10 N_WBL<10>_XI898/MM10_d N_WWLB<7>_XI898/MM10_g N_XI898/Q_XI898/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI898/MM11 N_WBLB<10>_XI898/MM11_d N_WWLB<7>_XI898/MM11_g
+ N_XI898/QB_XI898/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI898/MM1 N_XI898/Q_XI898/MM1_d N_XI898/QB_XI898/MM1_g N_GND_XI898/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI898/MM0 N_XI898/QB_XI898/MM0_d N_XI898/Q_XI898/MM0_g N_GND_XI898/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI898/MM9 N_XI898/NET08_XI898/MM9_d N_RWLB<7>_XI898/MM9_g N_RBL<10>_XI898/MM9_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI898/MM6 N_XI898/NET08_XI898/MM6_d N_XI898/QB_XI898/MM6_g N_VDD_XI898/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI898/MM5 N_XI898/Q_XI898/MM5_d N_XI898/QB_XI898/MM5_g N_VDD_XI898/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI898/MM4 N_XI898/QB_XI898/MM4_d N_XI898/Q_XI898/MM4_g N_VDD_XI898/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI897/MM8 N_XI897/NET08_XI897/MM8_d N_RWL<7>_XI897/MM8_g N_RBL<11>_XI897/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI897/MM7 N_XI897/NET08_XI897/MM7_d N_XI897/QB_XI897/MM7_g N_GND_XI897/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI897/MM10 N_WBL<11>_XI897/MM10_d N_WWLB<7>_XI897/MM10_g N_XI897/Q_XI897/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI897/MM11 N_WBLB<11>_XI897/MM11_d N_WWLB<7>_XI897/MM11_g
+ N_XI897/QB_XI897/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI897/MM1 N_XI897/Q_XI897/MM1_d N_XI897/QB_XI897/MM1_g N_GND_XI897/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI897/MM0 N_XI897/QB_XI897/MM0_d N_XI897/Q_XI897/MM0_g N_GND_XI897/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI897/MM9 N_XI897/NET08_XI897/MM9_d N_RWLB<7>_XI897/MM9_g N_RBL<11>_XI897/MM9_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI897/MM6 N_XI897/NET08_XI897/MM6_d N_XI897/QB_XI897/MM6_g N_VDD_XI897/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI897/MM5 N_XI897/Q_XI897/MM5_d N_XI897/QB_XI897/MM5_g N_VDD_XI897/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI897/MM4 N_XI897/QB_XI897/MM4_d N_XI897/Q_XI897/MM4_g N_VDD_XI897/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI896/MM8 N_XI896/NET08_XI896/MM8_d N_RWL<7>_XI896/MM8_g N_RBL<12>_XI896/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI896/MM7 N_XI896/NET08_XI896/MM7_d N_XI896/QB_XI896/MM7_g N_GND_XI896/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI896/MM10 N_WBL<12>_XI896/MM10_d N_WWLB<7>_XI896/MM10_g N_XI896/Q_XI896/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI896/MM11 N_WBLB<12>_XI896/MM11_d N_WWLB<7>_XI896/MM11_g
+ N_XI896/QB_XI896/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI896/MM1 N_XI896/Q_XI896/MM1_d N_XI896/QB_XI896/MM1_g N_GND_XI896/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI896/MM0 N_XI896/QB_XI896/MM0_d N_XI896/Q_XI896/MM0_g N_GND_XI896/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI896/MM9 N_XI896/NET08_XI896/MM9_d N_RWLB<7>_XI896/MM9_g N_RBL<12>_XI896/MM9_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI896/MM6 N_XI896/NET08_XI896/MM6_d N_XI896/QB_XI896/MM6_g N_VDD_XI896/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI896/MM5 N_XI896/Q_XI896/MM5_d N_XI896/QB_XI896/MM5_g N_VDD_XI896/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI896/MM4 N_XI896/QB_XI896/MM4_d N_XI896/Q_XI896/MM4_g N_VDD_XI896/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI885/MM8 N_XI885/NET08_XI885/MM8_d N_RWL<6>_XI885/MM8_g N_RBL<7>_XI885/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI885/MM7 N_XI885/NET08_XI885/MM7_d N_XI885/QB_XI885/MM7_g N_GND_XI885/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI885/MM10 N_WBL<7>_XI885/MM10_d N_WWLB<6>_XI885/MM10_g N_XI885/Q_XI885/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI885/MM11 N_WBLB<7>_XI885/MM11_d N_WWLB<6>_XI885/MM11_g
+ N_XI885/QB_XI885/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI885/MM1 N_XI885/Q_XI885/MM1_d N_XI885/QB_XI885/MM1_g N_GND_XI885/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI885/MM0 N_XI885/QB_XI885/MM0_d N_XI885/Q_XI885/MM0_g N_GND_XI885/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI885/MM9 N_XI885/NET08_XI885/MM9_d N_RWLB<6>_XI885/MM9_g N_RBL<7>_XI885/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI885/MM6 N_XI885/NET08_XI885/MM6_d N_XI885/QB_XI885/MM6_g N_VDD_XI885/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI885/MM5 N_XI885/Q_XI885/MM5_d N_XI885/QB_XI885/MM5_g N_VDD_XI885/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI885/MM4 N_XI885/QB_XI885/MM4_d N_XI885/Q_XI885/MM4_g N_VDD_XI885/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI884/MM8 N_XI884/NET08_XI884/MM8_d N_RWL<6>_XI884/MM8_g N_RBL<8>_XI884/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI884/MM7 N_XI884/NET08_XI884/MM7_d N_XI884/QB_XI884/MM7_g N_GND_XI884/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI884/MM10 N_WBL<8>_XI884/MM10_d N_WWLB<6>_XI884/MM10_g N_XI884/Q_XI884/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI884/MM11 N_WBLB<8>_XI884/MM11_d N_WWLB<6>_XI884/MM11_g
+ N_XI884/QB_XI884/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI884/MM1 N_XI884/Q_XI884/MM1_d N_XI884/QB_XI884/MM1_g N_GND_XI884/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI884/MM0 N_XI884/QB_XI884/MM0_d N_XI884/Q_XI884/MM0_g N_GND_XI884/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI884/MM9 N_XI884/NET08_XI884/MM9_d N_RWLB<6>_XI884/MM9_g N_RBL<8>_XI884/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI884/MM6 N_XI884/NET08_XI884/MM6_d N_XI884/QB_XI884/MM6_g N_VDD_XI884/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI884/MM5 N_XI884/Q_XI884/MM5_d N_XI884/QB_XI884/MM5_g N_VDD_XI884/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI884/MM4 N_XI884/QB_XI884/MM4_d N_XI884/Q_XI884/MM4_g N_VDD_XI884/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI883/MM8 N_XI883/NET08_XI883/MM8_d N_RWL<6>_XI883/MM8_g N_RBL<9>_XI883/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI883/MM7 N_XI883/NET08_XI883/MM7_d N_XI883/QB_XI883/MM7_g N_GND_XI883/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI883/MM10 N_WBL<9>_XI883/MM10_d N_WWLB<6>_XI883/MM10_g N_XI883/Q_XI883/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI883/MM11 N_WBLB<9>_XI883/MM11_d N_WWLB<6>_XI883/MM11_g
+ N_XI883/QB_XI883/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI883/MM1 N_XI883/Q_XI883/MM1_d N_XI883/QB_XI883/MM1_g N_GND_XI883/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI883/MM0 N_XI883/QB_XI883/MM0_d N_XI883/Q_XI883/MM0_g N_GND_XI883/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI883/MM9 N_XI883/NET08_XI883/MM9_d N_RWLB<6>_XI883/MM9_g N_RBL<9>_XI883/MM9_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI883/MM6 N_XI883/NET08_XI883/MM6_d N_XI883/QB_XI883/MM6_g N_VDD_XI883/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI883/MM5 N_XI883/Q_XI883/MM5_d N_XI883/QB_XI883/MM5_g N_VDD_XI883/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI883/MM4 N_XI883/QB_XI883/MM4_d N_XI883/Q_XI883/MM4_g N_VDD_XI883/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI882/MM8 N_XI882/NET08_XI882/MM8_d N_RWL<6>_XI882/MM8_g N_RBL<10>_XI882/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI882/MM7 N_XI882/NET08_XI882/MM7_d N_XI882/QB_XI882/MM7_g N_GND_XI882/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI882/MM10 N_WBL<10>_XI882/MM10_d N_WWLB<6>_XI882/MM10_g N_XI882/Q_XI882/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI882/MM11 N_WBLB<10>_XI882/MM11_d N_WWLB<6>_XI882/MM11_g
+ N_XI882/QB_XI882/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI882/MM1 N_XI882/Q_XI882/MM1_d N_XI882/QB_XI882/MM1_g N_GND_XI882/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI882/MM0 N_XI882/QB_XI882/MM0_d N_XI882/Q_XI882/MM0_g N_GND_XI882/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI882/MM9 N_XI882/NET08_XI882/MM9_d N_RWLB<6>_XI882/MM9_g N_RBL<10>_XI882/MM9_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI882/MM6 N_XI882/NET08_XI882/MM6_d N_XI882/QB_XI882/MM6_g N_VDD_XI882/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI882/MM5 N_XI882/Q_XI882/MM5_d N_XI882/QB_XI882/MM5_g N_VDD_XI882/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI882/MM4 N_XI882/QB_XI882/MM4_d N_XI882/Q_XI882/MM4_g N_VDD_XI882/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI919/MM8 N_XI919/NET08_XI919/MM8_d N_RWL<8>_XI919/MM8_g N_RBL<5>_XI919/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI919/MM7 N_XI919/NET08_XI919/MM7_d N_XI919/QB_XI919/MM7_g N_GND_XI919/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI919/MM10 N_WBL<5>_XI919/MM10_d N_WWLB<8>_XI919/MM10_g N_XI919/Q_XI919/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI919/MM11 N_WBLB<5>_XI919/MM11_d N_WWLB<8>_XI919/MM11_g
+ N_XI919/QB_XI919/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI919/MM1 N_XI919/Q_XI919/MM1_d N_XI919/QB_XI919/MM1_g N_GND_XI919/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI919/MM0 N_XI919/QB_XI919/MM0_d N_XI919/Q_XI919/MM0_g N_GND_XI919/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI919/MM9 N_XI919/NET08_XI919/MM9_d N_RWLB<8>_XI919/MM9_g N_RBL<5>_XI919/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI919/MM6 N_XI919/NET08_XI919/MM6_d N_XI919/QB_XI919/MM6_g N_VDD_XI919/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI919/MM5 N_XI919/Q_XI919/MM5_d N_XI919/QB_XI919/MM5_g N_VDD_XI919/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI919/MM4 N_XI919/QB_XI919/MM4_d N_XI919/Q_XI919/MM4_g N_VDD_XI919/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI918/MM8 N_XI918/NET08_XI918/MM8_d N_RWL<8>_XI918/MM8_g N_RBL<6>_XI918/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI918/MM7 N_XI918/NET08_XI918/MM7_d N_XI918/QB_XI918/MM7_g N_GND_XI918/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI918/MM10 N_WBL<6>_XI918/MM10_d N_WWLB<8>_XI918/MM10_g N_XI918/Q_XI918/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI918/MM11 N_WBLB<6>_XI918/MM11_d N_WWLB<8>_XI918/MM11_g
+ N_XI918/QB_XI918/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI918/MM1 N_XI918/Q_XI918/MM1_d N_XI918/QB_XI918/MM1_g N_GND_XI918/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI918/MM0 N_XI918/QB_XI918/MM0_d N_XI918/Q_XI918/MM0_g N_GND_XI918/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI918/MM9 N_XI918/NET08_XI918/MM9_d N_RWLB<8>_XI918/MM9_g N_RBL<6>_XI918/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI918/MM6 N_XI918/NET08_XI918/MM6_d N_XI918/QB_XI918/MM6_g N_VDD_XI918/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI918/MM5 N_XI918/Q_XI918/MM5_d N_XI918/QB_XI918/MM5_g N_VDD_XI918/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI918/MM4 N_XI918/QB_XI918/MM4_d N_XI918/Q_XI918/MM4_g N_VDD_XI918/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI917/MM8 N_XI917/NET08_XI917/MM8_d N_RWL<8>_XI917/MM8_g N_RBL<7>_XI917/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI917/MM7 N_XI917/NET08_XI917/MM7_d N_XI917/QB_XI917/MM7_g N_GND_XI917/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI917/MM10 N_WBL<7>_XI917/MM10_d N_WWLB<8>_XI917/MM10_g N_XI917/Q_XI917/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI917/MM11 N_WBLB<7>_XI917/MM11_d N_WWLB<8>_XI917/MM11_g
+ N_XI917/QB_XI917/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI917/MM1 N_XI917/Q_XI917/MM1_d N_XI917/QB_XI917/MM1_g N_GND_XI917/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI917/MM0 N_XI917/QB_XI917/MM0_d N_XI917/Q_XI917/MM0_g N_GND_XI917/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI917/MM9 N_XI917/NET08_XI917/MM9_d N_RWLB<8>_XI917/MM9_g N_RBL<7>_XI917/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI917/MM6 N_XI917/NET08_XI917/MM6_d N_XI917/QB_XI917/MM6_g N_VDD_XI917/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI917/MM5 N_XI917/Q_XI917/MM5_d N_XI917/QB_XI917/MM5_g N_VDD_XI917/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI917/MM4 N_XI917/QB_XI917/MM4_d N_XI917/Q_XI917/MM4_g N_VDD_XI917/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI916/MM8 N_XI916/NET08_XI916/MM8_d N_RWL<8>_XI916/MM8_g N_RBL<8>_XI916/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI916/MM7 N_XI916/NET08_XI916/MM7_d N_XI916/QB_XI916/MM7_g N_GND_XI916/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI916/MM10 N_WBL<8>_XI916/MM10_d N_WWLB<8>_XI916/MM10_g N_XI916/Q_XI916/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI916/MM11 N_WBLB<8>_XI916/MM11_d N_WWLB<8>_XI916/MM11_g
+ N_XI916/QB_XI916/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI916/MM1 N_XI916/Q_XI916/MM1_d N_XI916/QB_XI916/MM1_g N_GND_XI916/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI916/MM0 N_XI916/QB_XI916/MM0_d N_XI916/Q_XI916/MM0_g N_GND_XI916/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI916/MM9 N_XI916/NET08_XI916/MM9_d N_RWLB<8>_XI916/MM9_g N_RBL<8>_XI916/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI916/MM6 N_XI916/NET08_XI916/MM6_d N_XI916/QB_XI916/MM6_g N_VDD_XI916/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI916/MM5 N_XI916/Q_XI916/MM5_d N_XI916/QB_XI916/MM5_g N_VDD_XI916/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI916/MM4 N_XI916/QB_XI916/MM4_d N_XI916/Q_XI916/MM4_g N_VDD_XI916/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1028/MM8 N_XI1028/NET08_XI1028/MM8_d N_RWL<15>_XI1028/MM8_g
+ N_RBL<8>_XI1028/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1028/MM7 N_XI1028/NET08_XI1028/MM7_d N_XI1028/QB_XI1028/MM7_g
+ N_GND_XI1028/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1028/MM10 N_WBL<8>_XI1028/MM10_d N_WWLB<15>_XI1028/MM10_g
+ N_XI1028/Q_XI1028/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1028/MM11 N_WBLB<8>_XI1028/MM11_d N_WWLB<15>_XI1028/MM11_g
+ N_XI1028/QB_XI1028/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1028/MM1 N_XI1028/Q_XI1028/MM1_d N_XI1028/QB_XI1028/MM1_g N_GND_XI1028/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1028/MM0 N_XI1028/QB_XI1028/MM0_d N_XI1028/Q_XI1028/MM0_g N_GND_XI1028/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1028/MM9 N_XI1028/NET08_XI1028/MM9_d N_RWLB<15>_XI1028/MM9_g
+ N_RBL<8>_XI1028/MM9_s N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1028/MM6 N_XI1028/NET08_XI1028/MM6_d N_XI1028/QB_XI1028/MM6_g
+ N_VDD_XI1028/MM6_s N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1028/MM5 N_XI1028/Q_XI1028/MM5_d N_XI1028/QB_XI1028/MM5_g N_VDD_XI1028/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1028/MM4 N_XI1028/QB_XI1028/MM4_d N_XI1028/Q_XI1028/MM4_g N_VDD_XI1028/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI999/MM8 N_XI999/NET08_XI999/MM8_d N_RWL<13>_XI999/MM8_g N_RBL<5>_XI999/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI999/MM7 N_XI999/NET08_XI999/MM7_d N_XI999/QB_XI999/MM7_g N_GND_XI999/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI999/MM10 N_WBL<5>_XI999/MM10_d N_WWLB<13>_XI999/MM10_g N_XI999/Q_XI999/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI999/MM11 N_WBLB<5>_XI999/MM11_d N_WWLB<13>_XI999/MM11_g
+ N_XI999/QB_XI999/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI999/MM1 N_XI999/Q_XI999/MM1_d N_XI999/QB_XI999/MM1_g N_GND_XI999/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI999/MM0 N_XI999/QB_XI999/MM0_d N_XI999/Q_XI999/MM0_g N_GND_XI999/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI999/MM9 N_XI999/NET08_XI999/MM9_d N_RWLB<13>_XI999/MM9_g N_RBL<5>_XI999/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI999/MM6 N_XI999/NET08_XI999/MM6_d N_XI999/QB_XI999/MM6_g N_VDD_XI999/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI999/MM5 N_XI999/Q_XI999/MM5_d N_XI999/QB_XI999/MM5_g N_VDD_XI999/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI999/MM4 N_XI999/QB_XI999/MM4_d N_XI999/Q_XI999/MM4_g N_VDD_XI999/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI863/MM8 N_XI863/NET08_XI863/MM8_d N_RWL<5>_XI863/MM8_g N_RBL<13>_XI863/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI863/MM7 N_XI863/NET08_XI863/MM7_d N_XI863/QB_XI863/MM7_g N_GND_XI863/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI863/MM10 N_WBL<13>_XI863/MM10_d N_WWLB<5>_XI863/MM10_g N_XI863/Q_XI863/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI863/MM11 N_WBLB<13>_XI863/MM11_d N_WWLB<5>_XI863/MM11_g
+ N_XI863/QB_XI863/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI863/MM1 N_XI863/Q_XI863/MM1_d N_XI863/QB_XI863/MM1_g N_GND_XI863/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI863/MM0 N_XI863/QB_XI863/MM0_d N_XI863/Q_XI863/MM0_g N_GND_XI863/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI863/MM9 N_XI863/NET08_XI863/MM9_d N_RWLB<5>_XI863/MM9_g N_RBL<13>_XI863/MM9_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI863/MM6 N_XI863/NET08_XI863/MM6_d N_XI863/QB_XI863/MM6_g N_VDD_XI863/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI863/MM5 N_XI863/Q_XI863/MM5_d N_XI863/QB_XI863/MM5_g N_VDD_XI863/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI863/MM4 N_XI863/QB_XI863/MM4_d N_XI863/Q_XI863/MM4_g N_VDD_XI863/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI862/MM8 N_XI862/NET08_XI862/MM8_d N_RWL<5>_XI862/MM8_g N_RBL<14>_XI862/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI862/MM7 N_XI862/NET08_XI862/MM7_d N_XI862/QB_XI862/MM7_g N_GND_XI862/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI862/MM10 N_WBL<14>_XI862/MM10_d N_WWLB<5>_XI862/MM10_g N_XI862/Q_XI862/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI862/MM11 N_WBLB<14>_XI862/MM11_d N_WWLB<5>_XI862/MM11_g
+ N_XI862/QB_XI862/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI862/MM1 N_XI862/Q_XI862/MM1_d N_XI862/QB_XI862/MM1_g N_GND_XI862/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI862/MM0 N_XI862/QB_XI862/MM0_d N_XI862/Q_XI862/MM0_g N_GND_XI862/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI862/MM9 N_XI862/NET08_XI862/MM9_d N_RWLB<5>_XI862/MM9_g N_RBL<14>_XI862/MM9_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI862/MM6 N_XI862/NET08_XI862/MM6_d N_XI862/QB_XI862/MM6_g N_VDD_XI862/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI862/MM5 N_XI862/Q_XI862/MM5_d N_XI862/QB_XI862/MM5_g N_VDD_XI862/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI862/MM4 N_XI862/QB_XI862/MM4_d N_XI862/Q_XI862/MM4_g N_VDD_XI862/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI861/MM8 N_XI861/NET08_XI861/MM8_d N_RWL<4>_XI861/MM8_g N_RBL<15>_XI861/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI861/MM7 N_XI861/NET08_XI861/MM7_d N_XI861/QB_XI861/MM7_g N_GND_XI861/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI861/MM10 N_WBL<15>_XI861/MM10_d N_WWLB<4>_XI861/MM10_g N_XI861/Q_XI861/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI861/MM11 N_WBLB<15>_XI861/MM11_d N_WWLB<4>_XI861/MM11_g
+ N_XI861/QB_XI861/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI861/MM1 N_XI861/Q_XI861/MM1_d N_XI861/QB_XI861/MM1_g N_GND_XI861/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI861/MM0 N_XI861/QB_XI861/MM0_d N_XI861/Q_XI861/MM0_g N_GND_XI861/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI861/MM9 N_XI861/NET08_XI861/MM9_d N_RWLB<4>_XI861/MM9_g N_RBL<15>_XI861/MM9_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI861/MM6 N_XI861/NET08_XI861/MM6_d N_XI861/QB_XI861/MM6_g N_VDD_XI861/MM6_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI861/MM5 N_XI861/Q_XI861/MM5_d N_XI861/QB_XI861/MM5_g N_VDD_XI861/MM5_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI861/MM4 N_XI861/QB_XI861/MM4_d N_XI861/Q_XI861/MM4_g N_VDD_XI861/MM4_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI860/MM8 N_XI860/NET08_XI860/MM8_d N_RWL<4>_XI860/MM8_g N_RBL<0>_XI860/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI860/MM7 N_XI860/NET08_XI860/MM7_d N_XI860/QB_XI860/MM7_g N_GND_XI860/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI860/MM10 N_WBL<0>_XI860/MM10_d N_WWLB<4>_XI860/MM10_g N_XI860/Q_XI860/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI860/MM11 N_WBLB<0>_XI860/MM11_d N_WWLB<4>_XI860/MM11_g
+ N_XI860/QB_XI860/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI860/MM1 N_XI860/Q_XI860/MM1_d N_XI860/QB_XI860/MM1_g N_GND_XI860/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI860/MM0 N_XI860/QB_XI860/MM0_d N_XI860/Q_XI860/MM0_g N_GND_XI860/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI860/MM9 N_XI860/NET08_XI860/MM9_d N_RWLB<4>_XI860/MM9_g N_RBL<0>_XI860/MM9_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI860/MM6 N_XI860/NET08_XI860/MM6_d N_XI860/QB_XI860/MM6_g N_VDD_XI860/MM6_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI860/MM5 N_XI860/Q_XI860/MM5_d N_XI860/QB_XI860/MM5_g N_VDD_XI860/MM5_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI860/MM4 N_XI860/QB_XI860/MM4_d N_XI860/Q_XI860/MM4_g N_VDD_XI860/MM4_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI893/MM8 N_XI893/NET08_XI893/MM8_d N_RWL<6>_XI893/MM8_g N_RBL<15>_XI893/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI893/MM7 N_XI893/NET08_XI893/MM7_d N_XI893/QB_XI893/MM7_g N_GND_XI893/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI893/MM10 N_WBL<15>_XI893/MM10_d N_WWLB<6>_XI893/MM10_g N_XI893/Q_XI893/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI893/MM11 N_WBLB<15>_XI893/MM11_d N_WWLB<6>_XI893/MM11_g
+ N_XI893/QB_XI893/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI893/MM1 N_XI893/Q_XI893/MM1_d N_XI893/QB_XI893/MM1_g N_GND_XI893/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI893/MM0 N_XI893/QB_XI893/MM0_d N_XI893/Q_XI893/MM0_g N_GND_XI893/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI893/MM9 N_XI893/NET08_XI893/MM9_d N_RWLB<6>_XI893/MM9_g N_RBL<15>_XI893/MM9_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI893/MM6 N_XI893/NET08_XI893/MM6_d N_XI893/QB_XI893/MM6_g N_VDD_XI893/MM6_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI893/MM5 N_XI893/Q_XI893/MM5_d N_XI893/QB_XI893/MM5_g N_VDD_XI893/MM5_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI893/MM4 N_XI893/QB_XI893/MM4_d N_XI893/Q_XI893/MM4_g N_VDD_XI893/MM4_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI892/MM8 N_XI892/NET08_XI892/MM8_d N_RWL<6>_XI892/MM8_g N_RBL<0>_XI892/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI892/MM7 N_XI892/NET08_XI892/MM7_d N_XI892/QB_XI892/MM7_g N_GND_XI892/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI892/MM10 N_WBL<0>_XI892/MM10_d N_WWLB<6>_XI892/MM10_g N_XI892/Q_XI892/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI892/MM11 N_WBLB<0>_XI892/MM11_d N_WWLB<6>_XI892/MM11_g
+ N_XI892/QB_XI892/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI892/MM1 N_XI892/Q_XI892/MM1_d N_XI892/QB_XI892/MM1_g N_GND_XI892/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI892/MM0 N_XI892/QB_XI892/MM0_d N_XI892/Q_XI892/MM0_g N_GND_XI892/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI892/MM9 N_XI892/NET08_XI892/MM9_d N_RWLB<6>_XI892/MM9_g N_RBL<0>_XI892/MM9_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI892/MM6 N_XI892/NET08_XI892/MM6_d N_XI892/QB_XI892/MM6_g N_VDD_XI892/MM6_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI892/MM5 N_XI892/Q_XI892/MM5_d N_XI892/QB_XI892/MM5_g N_VDD_XI892/MM5_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI892/MM4 N_XI892/QB_XI892/MM4_d N_XI892/Q_XI892/MM4_g N_VDD_XI892/MM4_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI891/MM8 N_XI891/NET08_XI891/MM8_d N_RWL<6>_XI891/MM8_g N_RBL<1>_XI891/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI891/MM7 N_XI891/NET08_XI891/MM7_d N_XI891/QB_XI891/MM7_g N_GND_XI891/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI891/MM10 N_WBL<1>_XI891/MM10_d N_WWLB<6>_XI891/MM10_g N_XI891/Q_XI891/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI891/MM11 N_WBLB<1>_XI891/MM11_d N_WWLB<6>_XI891/MM11_g
+ N_XI891/QB_XI891/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI891/MM1 N_XI891/Q_XI891/MM1_d N_XI891/QB_XI891/MM1_g N_GND_XI891/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI891/MM0 N_XI891/QB_XI891/MM0_d N_XI891/Q_XI891/MM0_g N_GND_XI891/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI891/MM9 N_XI891/NET08_XI891/MM9_d N_RWLB<6>_XI891/MM9_g N_RBL<1>_XI891/MM9_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI891/MM6 N_XI891/NET08_XI891/MM6_d N_XI891/QB_XI891/MM6_g N_VDD_XI891/MM6_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI891/MM5 N_XI891/Q_XI891/MM5_d N_XI891/QB_XI891/MM5_g N_VDD_XI891/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI891/MM4 N_XI891/QB_XI891/MM4_d N_XI891/Q_XI891/MM4_g N_VDD_XI891/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI879/MM8 N_XI879/NET08_XI879/MM8_d N_RWL<6>_XI879/MM8_g N_RBL<13>_XI879/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI879/MM7 N_XI879/NET08_XI879/MM7_d N_XI879/QB_XI879/MM7_g N_GND_XI879/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI879/MM10 N_WBL<13>_XI879/MM10_d N_WWLB<6>_XI879/MM10_g N_XI879/Q_XI879/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI879/MM11 N_WBLB<13>_XI879/MM11_d N_WWLB<6>_XI879/MM11_g
+ N_XI879/QB_XI879/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI879/MM1 N_XI879/Q_XI879/MM1_d N_XI879/QB_XI879/MM1_g N_GND_XI879/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI879/MM0 N_XI879/QB_XI879/MM0_d N_XI879/Q_XI879/MM0_g N_GND_XI879/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI879/MM9 N_XI879/NET08_XI879/MM9_d N_RWLB<6>_XI879/MM9_g N_RBL<13>_XI879/MM9_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI879/MM6 N_XI879/NET08_XI879/MM6_d N_XI879/QB_XI879/MM6_g N_VDD_XI879/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI879/MM5 N_XI879/Q_XI879/MM5_d N_XI879/QB_XI879/MM5_g N_VDD_XI879/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI879/MM4 N_XI879/QB_XI879/MM4_d N_XI879/Q_XI879/MM4_g N_VDD_XI879/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI878/MM8 N_XI878/NET08_XI878/MM8_d N_RWL<6>_XI878/MM8_g N_RBL<14>_XI878/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI878/MM7 N_XI878/NET08_XI878/MM7_d N_XI878/QB_XI878/MM7_g N_GND_XI878/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI878/MM10 N_WBL<14>_XI878/MM10_d N_WWLB<6>_XI878/MM10_g N_XI878/Q_XI878/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI878/MM11 N_WBLB<14>_XI878/MM11_d N_WWLB<6>_XI878/MM11_g
+ N_XI878/QB_XI878/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI878/MM1 N_XI878/Q_XI878/MM1_d N_XI878/QB_XI878/MM1_g N_GND_XI878/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI878/MM0 N_XI878/QB_XI878/MM0_d N_XI878/Q_XI878/MM0_g N_GND_XI878/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI878/MM9 N_XI878/NET08_XI878/MM9_d N_RWLB<6>_XI878/MM9_g N_RBL<14>_XI878/MM9_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI878/MM6 N_XI878/NET08_XI878/MM6_d N_XI878/QB_XI878/MM6_g N_VDD_XI878/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI878/MM5 N_XI878/Q_XI878/MM5_d N_XI878/QB_XI878/MM5_g N_VDD_XI878/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI878/MM4 N_XI878/QB_XI878/MM4_d N_XI878/Q_XI878/MM4_g N_VDD_XI878/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI877/MM8 N_XI877/NET08_XI877/MM8_d N_RWL<5>_XI877/MM8_g N_RBL<15>_XI877/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI877/MM7 N_XI877/NET08_XI877/MM7_d N_XI877/QB_XI877/MM7_g N_GND_XI877/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI877/MM10 N_WBL<15>_XI877/MM10_d N_WWLB<5>_XI877/MM10_g N_XI877/Q_XI877/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI877/MM11 N_WBLB<15>_XI877/MM11_d N_WWLB<5>_XI877/MM11_g
+ N_XI877/QB_XI877/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI877/MM1 N_XI877/Q_XI877/MM1_d N_XI877/QB_XI877/MM1_g N_GND_XI877/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI877/MM0 N_XI877/QB_XI877/MM0_d N_XI877/Q_XI877/MM0_g N_GND_XI877/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI877/MM9 N_XI877/NET08_XI877/MM9_d N_RWLB<5>_XI877/MM9_g N_RBL<15>_XI877/MM9_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI877/MM6 N_XI877/NET08_XI877/MM6_d N_XI877/QB_XI877/MM6_g N_VDD_XI877/MM6_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI877/MM5 N_XI877/Q_XI877/MM5_d N_XI877/QB_XI877/MM5_g N_VDD_XI877/MM5_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI877/MM4 N_XI877/QB_XI877/MM4_d N_XI877/Q_XI877/MM4_g N_VDD_XI877/MM4_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI876/MM8 N_XI876/NET08_XI876/MM8_d N_RWL<5>_XI876/MM8_g N_RBL<0>_XI876/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI876/MM7 N_XI876/NET08_XI876/MM7_d N_XI876/QB_XI876/MM7_g N_GND_XI876/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI876/MM10 N_WBL<0>_XI876/MM10_d N_WWLB<5>_XI876/MM10_g N_XI876/Q_XI876/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI876/MM11 N_WBLB<0>_XI876/MM11_d N_WWLB<5>_XI876/MM11_g
+ N_XI876/QB_XI876/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI876/MM1 N_XI876/Q_XI876/MM1_d N_XI876/QB_XI876/MM1_g N_GND_XI876/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI876/MM0 N_XI876/QB_XI876/MM0_d N_XI876/Q_XI876/MM0_g N_GND_XI876/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI876/MM9 N_XI876/NET08_XI876/MM9_d N_RWLB<5>_XI876/MM9_g N_RBL<0>_XI876/MM9_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI876/MM6 N_XI876/NET08_XI876/MM6_d N_XI876/QB_XI876/MM6_g N_VDD_XI876/MM6_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI876/MM5 N_XI876/Q_XI876/MM5_d N_XI876/QB_XI876/MM5_g N_VDD_XI876/MM5_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI876/MM4 N_XI876/QB_XI876/MM4_d N_XI876/Q_XI876/MM4_g N_VDD_XI876/MM4_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI881/MM8 N_XI881/NET08_XI881/MM8_d N_RWL<6>_XI881/MM8_g N_RBL<11>_XI881/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI881/MM7 N_XI881/NET08_XI881/MM7_d N_XI881/QB_XI881/MM7_g N_GND_XI881/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI881/MM10 N_WBL<11>_XI881/MM10_d N_WWLB<6>_XI881/MM10_g N_XI881/Q_XI881/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI881/MM11 N_WBLB<11>_XI881/MM11_d N_WWLB<6>_XI881/MM11_g
+ N_XI881/QB_XI881/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI881/MM1 N_XI881/Q_XI881/MM1_d N_XI881/QB_XI881/MM1_g N_GND_XI881/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI881/MM0 N_XI881/QB_XI881/MM0_d N_XI881/Q_XI881/MM0_g N_GND_XI881/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI881/MM9 N_XI881/NET08_XI881/MM9_d N_RWLB<6>_XI881/MM9_g N_RBL<11>_XI881/MM9_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI881/MM6 N_XI881/NET08_XI881/MM6_d N_XI881/QB_XI881/MM6_g N_VDD_XI881/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI881/MM5 N_XI881/Q_XI881/MM5_d N_XI881/QB_XI881/MM5_g N_VDD_XI881/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI881/MM4 N_XI881/QB_XI881/MM4_d N_XI881/Q_XI881/MM4_g N_VDD_XI881/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI915/MM8 N_XI915/NET08_XI915/MM8_d N_RWL<8>_XI915/MM8_g N_RBL<9>_XI915/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI915/MM7 N_XI915/NET08_XI915/MM7_d N_XI915/QB_XI915/MM7_g N_GND_XI915/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI915/MM10 N_WBL<9>_XI915/MM10_d N_WWLB<8>_XI915/MM10_g N_XI915/Q_XI915/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI915/MM11 N_WBLB<9>_XI915/MM11_d N_WWLB<8>_XI915/MM11_g
+ N_XI915/QB_XI915/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI915/MM1 N_XI915/Q_XI915/MM1_d N_XI915/QB_XI915/MM1_g N_GND_XI915/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI915/MM0 N_XI915/QB_XI915/MM0_d N_XI915/Q_XI915/MM0_g N_GND_XI915/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI915/MM9 N_XI915/NET08_XI915/MM9_d N_RWLB<8>_XI915/MM9_g N_RBL<9>_XI915/MM9_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI915/MM6 N_XI915/NET08_XI915/MM6_d N_XI915/QB_XI915/MM6_g N_VDD_XI915/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI915/MM5 N_XI915/Q_XI915/MM5_d N_XI915/QB_XI915/MM5_g N_VDD_XI915/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI915/MM4 N_XI915/QB_XI915/MM4_d N_XI915/Q_XI915/MM4_g N_VDD_XI915/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI914/MM8 N_XI914/NET08_XI914/MM8_d N_RWL<8>_XI914/MM8_g N_RBL<10>_XI914/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI914/MM7 N_XI914/NET08_XI914/MM7_d N_XI914/QB_XI914/MM7_g N_GND_XI914/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI914/MM10 N_WBL<10>_XI914/MM10_d N_WWLB<8>_XI914/MM10_g N_XI914/Q_XI914/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI914/MM11 N_WBLB<10>_XI914/MM11_d N_WWLB<8>_XI914/MM11_g
+ N_XI914/QB_XI914/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI914/MM1 N_XI914/Q_XI914/MM1_d N_XI914/QB_XI914/MM1_g N_GND_XI914/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI914/MM0 N_XI914/QB_XI914/MM0_d N_XI914/Q_XI914/MM0_g N_GND_XI914/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI914/MM9 N_XI914/NET08_XI914/MM9_d N_RWLB<8>_XI914/MM9_g N_RBL<10>_XI914/MM9_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI914/MM6 N_XI914/NET08_XI914/MM6_d N_XI914/QB_XI914/MM6_g N_VDD_XI914/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI914/MM5 N_XI914/Q_XI914/MM5_d N_XI914/QB_XI914/MM5_g N_VDD_XI914/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI914/MM4 N_XI914/QB_XI914/MM4_d N_XI914/Q_XI914/MM4_g N_VDD_XI914/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI913/MM8 N_XI913/NET08_XI913/MM8_d N_RWL<8>_XI913/MM8_g N_RBL<11>_XI913/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI913/MM7 N_XI913/NET08_XI913/MM7_d N_XI913/QB_XI913/MM7_g N_GND_XI913/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI913/MM10 N_WBL<11>_XI913/MM10_d N_WWLB<8>_XI913/MM10_g N_XI913/Q_XI913/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI913/MM11 N_WBLB<11>_XI913/MM11_d N_WWLB<8>_XI913/MM11_g
+ N_XI913/QB_XI913/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI913/MM1 N_XI913/Q_XI913/MM1_d N_XI913/QB_XI913/MM1_g N_GND_XI913/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI913/MM0 N_XI913/QB_XI913/MM0_d N_XI913/Q_XI913/MM0_g N_GND_XI913/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI913/MM9 N_XI913/NET08_XI913/MM9_d N_RWLB<8>_XI913/MM9_g N_RBL<11>_XI913/MM9_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI913/MM6 N_XI913/NET08_XI913/MM6_d N_XI913/QB_XI913/MM6_g N_VDD_XI913/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI913/MM5 N_XI913/Q_XI913/MM5_d N_XI913/QB_XI913/MM5_g N_VDD_XI913/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI913/MM4 N_XI913/QB_XI913/MM4_d N_XI913/Q_XI913/MM4_g N_VDD_XI913/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI912/MM8 N_XI912/NET08_XI912/MM8_d N_RWL<8>_XI912/MM8_g N_RBL<12>_XI912/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI912/MM7 N_XI912/NET08_XI912/MM7_d N_XI912/QB_XI912/MM7_g N_GND_XI912/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI912/MM10 N_WBL<12>_XI912/MM10_d N_WWLB<8>_XI912/MM10_g N_XI912/Q_XI912/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI912/MM11 N_WBLB<12>_XI912/MM11_d N_WWLB<8>_XI912/MM11_g
+ N_XI912/QB_XI912/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI912/MM1 N_XI912/Q_XI912/MM1_d N_XI912/QB_XI912/MM1_g N_GND_XI912/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI912/MM0 N_XI912/QB_XI912/MM0_d N_XI912/Q_XI912/MM0_g N_GND_XI912/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI912/MM9 N_XI912/NET08_XI912/MM9_d N_RWLB<8>_XI912/MM9_g N_RBL<12>_XI912/MM9_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI912/MM6 N_XI912/NET08_XI912/MM6_d N_XI912/QB_XI912/MM6_g N_VDD_XI912/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI912/MM5 N_XI912/Q_XI912/MM5_d N_XI912/QB_XI912/MM5_g N_VDD_XI912/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI912/MM4 N_XI912/QB_XI912/MM4_d N_XI912/Q_XI912/MM4_g N_VDD_XI912/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1027/MM8 N_XI1027/NET08_XI1027/MM8_d N_RWL<15>_XI1027/MM8_g
+ N_RBL<9>_XI1027/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1027/MM7 N_XI1027/NET08_XI1027/MM7_d N_XI1027/QB_XI1027/MM7_g
+ N_GND_XI1027/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1027/MM10 N_WBL<9>_XI1027/MM10_d N_WWLB<15>_XI1027/MM10_g
+ N_XI1027/Q_XI1027/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1027/MM11 N_WBLB<9>_XI1027/MM11_d N_WWLB<15>_XI1027/MM11_g
+ N_XI1027/QB_XI1027/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1027/MM1 N_XI1027/Q_XI1027/MM1_d N_XI1027/QB_XI1027/MM1_g N_GND_XI1027/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1027/MM0 N_XI1027/QB_XI1027/MM0_d N_XI1027/Q_XI1027/MM0_g N_GND_XI1027/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1027/MM9 N_XI1027/NET08_XI1027/MM9_d N_RWLB<15>_XI1027/MM9_g
+ N_RBL<9>_XI1027/MM9_s N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1027/MM6 N_XI1027/NET08_XI1027/MM6_d N_XI1027/QB_XI1027/MM6_g
+ N_VDD_XI1027/MM6_s N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1027/MM5 N_XI1027/Q_XI1027/MM5_d N_XI1027/QB_XI1027/MM5_g N_VDD_XI1027/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1027/MM4 N_XI1027/QB_XI1027/MM4_d N_XI1027/Q_XI1027/MM4_g N_VDD_XI1027/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1000/MM8 N_XI1000/NET08_XI1000/MM8_d N_RWL<13>_XI1000/MM8_g
+ N_RBL<4>_XI1000/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1000/MM7 N_XI1000/NET08_XI1000/MM7_d N_XI1000/QB_XI1000/MM7_g
+ N_GND_XI1000/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1000/MM10 N_WBL<4>_XI1000/MM10_d N_WWLB<13>_XI1000/MM10_g
+ N_XI1000/Q_XI1000/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1000/MM11 N_WBLB<4>_XI1000/MM11_d N_WWLB<13>_XI1000/MM11_g
+ N_XI1000/QB_XI1000/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1000/MM1 N_XI1000/Q_XI1000/MM1_d N_XI1000/QB_XI1000/MM1_g N_GND_XI1000/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1000/MM0 N_XI1000/QB_XI1000/MM0_d N_XI1000/Q_XI1000/MM0_g N_GND_XI1000/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1000/MM9 N_XI1000/NET08_XI1000/MM9_d N_RWLB<13>_XI1000/MM9_g
+ N_RBL<4>_XI1000/MM9_s N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1000/MM6 N_XI1000/NET08_XI1000/MM6_d N_XI1000/QB_XI1000/MM6_g
+ N_VDD_XI1000/MM6_s N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1000/MM5 N_XI1000/Q_XI1000/MM5_d N_XI1000/QB_XI1000/MM5_g N_VDD_XI1000/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1000/MM4 N_XI1000/QB_XI1000/MM4_d N_XI1000/Q_XI1000/MM4_g N_VDD_XI1000/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI859/MM8 N_XI859/NET08_XI859/MM8_d N_RWL<4>_XI859/MM8_g N_RBL<1>_XI859/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI859/MM7 N_XI859/NET08_XI859/MM7_d N_XI859/QB_XI859/MM7_g N_GND_XI859/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI859/MM10 N_WBL<1>_XI859/MM10_d N_WWLB<4>_XI859/MM10_g N_XI859/Q_XI859/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI859/MM11 N_WBLB<1>_XI859/MM11_d N_WWLB<4>_XI859/MM11_g
+ N_XI859/QB_XI859/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI859/MM1 N_XI859/Q_XI859/MM1_d N_XI859/QB_XI859/MM1_g N_GND_XI859/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI859/MM0 N_XI859/QB_XI859/MM0_d N_XI859/Q_XI859/MM0_g N_GND_XI859/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI859/MM9 N_XI859/NET08_XI859/MM9_d N_RWLB<4>_XI859/MM9_g N_RBL<1>_XI859/MM9_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI859/MM6 N_XI859/NET08_XI859/MM6_d N_XI859/QB_XI859/MM6_g N_VDD_XI859/MM6_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI859/MM5 N_XI859/Q_XI859/MM5_d N_XI859/QB_XI859/MM5_g N_VDD_XI859/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI859/MM4 N_XI859/QB_XI859/MM4_d N_XI859/Q_XI859/MM4_g N_VDD_XI859/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI858/MM8 N_XI858/NET08_XI858/MM8_d N_RWL<4>_XI858/MM8_g N_RBL<2>_XI858/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI858/MM7 N_XI858/NET08_XI858/MM7_d N_XI858/QB_XI858/MM7_g N_GND_XI858/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI858/MM10 N_WBL<2>_XI858/MM10_d N_WWLB<4>_XI858/MM10_g N_XI858/Q_XI858/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI858/MM11 N_WBLB<2>_XI858/MM11_d N_WWLB<4>_XI858/MM11_g
+ N_XI858/QB_XI858/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI858/MM1 N_XI858/Q_XI858/MM1_d N_XI858/QB_XI858/MM1_g N_GND_XI858/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI858/MM0 N_XI858/QB_XI858/MM0_d N_XI858/Q_XI858/MM0_g N_GND_XI858/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI858/MM9 N_XI858/NET08_XI858/MM9_d N_RWLB<4>_XI858/MM9_g N_RBL<2>_XI858/MM9_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI858/MM6 N_XI858/NET08_XI858/MM6_d N_XI858/QB_XI858/MM6_g N_VDD_XI858/MM6_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI858/MM5 N_XI858/Q_XI858/MM5_d N_XI858/QB_XI858/MM5_g N_VDD_XI858/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI858/MM4 N_XI858/QB_XI858/MM4_d N_XI858/Q_XI858/MM4_g N_VDD_XI858/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI857/MM8 N_XI857/NET08_XI857/MM8_d N_RWL<4>_XI857/MM8_g N_RBL<3>_XI857/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI857/MM7 N_XI857/NET08_XI857/MM7_d N_XI857/QB_XI857/MM7_g N_GND_XI857/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI857/MM10 N_WBL<3>_XI857/MM10_d N_WWLB<4>_XI857/MM10_g N_XI857/Q_XI857/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI857/MM11 N_WBLB<3>_XI857/MM11_d N_WWLB<4>_XI857/MM11_g
+ N_XI857/QB_XI857/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI857/MM1 N_XI857/Q_XI857/MM1_d N_XI857/QB_XI857/MM1_g N_GND_XI857/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI857/MM0 N_XI857/QB_XI857/MM0_d N_XI857/Q_XI857/MM0_g N_GND_XI857/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI857/MM9 N_XI857/NET08_XI857/MM9_d N_RWLB<4>_XI857/MM9_g N_RBL<3>_XI857/MM9_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI857/MM6 N_XI857/NET08_XI857/MM6_d N_XI857/QB_XI857/MM6_g N_VDD_XI857/MM6_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI857/MM5 N_XI857/Q_XI857/MM5_d N_XI857/QB_XI857/MM5_g N_VDD_XI857/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI857/MM4 N_XI857/QB_XI857/MM4_d N_XI857/Q_XI857/MM4_g N_VDD_XI857/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI856/MM8 N_XI856/NET08_XI856/MM8_d N_RWL<4>_XI856/MM8_g N_RBL<4>_XI856/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI856/MM7 N_XI856/NET08_XI856/MM7_d N_XI856/QB_XI856/MM7_g N_GND_XI856/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI856/MM10 N_WBL<4>_XI856/MM10_d N_WWLB<4>_XI856/MM10_g N_XI856/Q_XI856/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI856/MM11 N_WBLB<4>_XI856/MM11_d N_WWLB<4>_XI856/MM11_g
+ N_XI856/QB_XI856/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI856/MM1 N_XI856/Q_XI856/MM1_d N_XI856/QB_XI856/MM1_g N_GND_XI856/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI856/MM0 N_XI856/QB_XI856/MM0_d N_XI856/Q_XI856/MM0_g N_GND_XI856/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI856/MM9 N_XI856/NET08_XI856/MM9_d N_RWLB<4>_XI856/MM9_g N_RBL<4>_XI856/MM9_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI856/MM6 N_XI856/NET08_XI856/MM6_d N_XI856/QB_XI856/MM6_g N_VDD_XI856/MM6_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI856/MM5 N_XI856/Q_XI856/MM5_d N_XI856/QB_XI856/MM5_g N_VDD_XI856/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI856/MM4 N_XI856/QB_XI856/MM4_d N_XI856/Q_XI856/MM4_g N_VDD_XI856/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI887/MM8 N_XI887/NET08_XI887/MM8_d N_RWL<6>_XI887/MM8_g N_RBL<5>_XI887/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI887/MM7 N_XI887/NET08_XI887/MM7_d N_XI887/QB_XI887/MM7_g N_GND_XI887/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI887/MM10 N_WBL<5>_XI887/MM10_d N_WWLB<6>_XI887/MM10_g N_XI887/Q_XI887/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI887/MM11 N_WBLB<5>_XI887/MM11_d N_WWLB<6>_XI887/MM11_g
+ N_XI887/QB_XI887/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI887/MM1 N_XI887/Q_XI887/MM1_d N_XI887/QB_XI887/MM1_g N_GND_XI887/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI887/MM0 N_XI887/QB_XI887/MM0_d N_XI887/Q_XI887/MM0_g N_GND_XI887/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI887/MM9 N_XI887/NET08_XI887/MM9_d N_RWLB<6>_XI887/MM9_g N_RBL<5>_XI887/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI887/MM6 N_XI887/NET08_XI887/MM6_d N_XI887/QB_XI887/MM6_g N_VDD_XI887/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI887/MM5 N_XI887/Q_XI887/MM5_d N_XI887/QB_XI887/MM5_g N_VDD_XI887/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI887/MM4 N_XI887/QB_XI887/MM4_d N_XI887/Q_XI887/MM4_g N_VDD_XI887/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI886/MM8 N_XI886/NET08_XI886/MM8_d N_RWL<6>_XI886/MM8_g N_RBL<6>_XI886/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI886/MM7 N_XI886/NET08_XI886/MM7_d N_XI886/QB_XI886/MM7_g N_GND_XI886/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI886/MM10 N_WBL<6>_XI886/MM10_d N_WWLB<6>_XI886/MM10_g N_XI886/Q_XI886/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI886/MM11 N_WBLB<6>_XI886/MM11_d N_WWLB<6>_XI886/MM11_g
+ N_XI886/QB_XI886/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI886/MM1 N_XI886/Q_XI886/MM1_d N_XI886/QB_XI886/MM1_g N_GND_XI886/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI886/MM0 N_XI886/QB_XI886/MM0_d N_XI886/Q_XI886/MM0_g N_GND_XI886/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI886/MM9 N_XI886/NET08_XI886/MM9_d N_RWLB<6>_XI886/MM9_g N_RBL<6>_XI886/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI886/MM6 N_XI886/NET08_XI886/MM6_d N_XI886/QB_XI886/MM6_g N_VDD_XI886/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI886/MM5 N_XI886/Q_XI886/MM5_d N_XI886/QB_XI886/MM5_g N_VDD_XI886/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI886/MM4 N_XI886/QB_XI886/MM4_d N_XI886/Q_XI886/MM4_g N_VDD_XI886/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI831/MM8 N_XI831/NET08_XI831/MM8_d N_RWL<3>_XI831/MM8_g N_RBL<13>_XI831/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI831/MM7 N_XI831/NET08_XI831/MM7_d N_XI831/QB_XI831/MM7_g N_GND_XI831/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI831/MM10 N_WBL<13>_XI831/MM10_d N_WWLB<3>_XI831/MM10_g N_XI831/Q_XI831/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI831/MM11 N_WBLB<13>_XI831/MM11_d N_WWLB<3>_XI831/MM11_g
+ N_XI831/QB_XI831/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI831/MM1 N_XI831/Q_XI831/MM1_d N_XI831/QB_XI831/MM1_g N_GND_XI831/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI831/MM0 N_XI831/QB_XI831/MM0_d N_XI831/Q_XI831/MM0_g N_GND_XI831/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI831/MM9 N_XI831/NET08_XI831/MM9_d N_RWLB<3>_XI831/MM9_g N_RBL<13>_XI831/MM9_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI831/MM6 N_XI831/NET08_XI831/MM6_d N_XI831/QB_XI831/MM6_g N_VDD_XI831/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI831/MM5 N_XI831/Q_XI831/MM5_d N_XI831/QB_XI831/MM5_g N_VDD_XI831/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI831/MM4 N_XI831/QB_XI831/MM4_d N_XI831/Q_XI831/MM4_g N_VDD_XI831/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI830/MM8 N_XI830/NET08_XI830/MM8_d N_RWL<3>_XI830/MM8_g N_RBL<14>_XI830/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI830/MM7 N_XI830/NET08_XI830/MM7_d N_XI830/QB_XI830/MM7_g N_GND_XI830/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI830/MM10 N_WBL<14>_XI830/MM10_d N_WWLB<3>_XI830/MM10_g N_XI830/Q_XI830/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI830/MM11 N_WBLB<14>_XI830/MM11_d N_WWLB<3>_XI830/MM11_g
+ N_XI830/QB_XI830/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI830/MM1 N_XI830/Q_XI830/MM1_d N_XI830/QB_XI830/MM1_g N_GND_XI830/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI830/MM0 N_XI830/QB_XI830/MM0_d N_XI830/Q_XI830/MM0_g N_GND_XI830/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI830/MM9 N_XI830/NET08_XI830/MM9_d N_RWLB<3>_XI830/MM9_g N_RBL<14>_XI830/MM9_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI830/MM6 N_XI830/NET08_XI830/MM6_d N_XI830/QB_XI830/MM6_g N_VDD_XI830/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI830/MM5 N_XI830/Q_XI830/MM5_d N_XI830/QB_XI830/MM5_g N_VDD_XI830/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI830/MM4 N_XI830/QB_XI830/MM4_d N_XI830/Q_XI830/MM4_g N_VDD_XI830/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI829/MM8 N_XI829/NET08_XI829/MM8_d N_RWL<2>_XI829/MM8_g N_RBL<15>_XI829/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI829/MM7 N_XI829/NET08_XI829/MM7_d N_XI829/QB_XI829/MM7_g N_GND_XI829/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI829/MM10 N_WBL<15>_XI829/MM10_d N_WWLB<2>_XI829/MM10_g N_XI829/Q_XI829/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI829/MM11 N_WBLB<15>_XI829/MM11_d N_WWLB<2>_XI829/MM11_g
+ N_XI829/QB_XI829/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI829/MM1 N_XI829/Q_XI829/MM1_d N_XI829/QB_XI829/MM1_g N_GND_XI829/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI829/MM0 N_XI829/QB_XI829/MM0_d N_XI829/Q_XI829/MM0_g N_GND_XI829/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI829/MM9 N_XI829/NET08_XI829/MM9_d N_RWLB<2>_XI829/MM9_g N_RBL<15>_XI829/MM9_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI829/MM6 N_XI829/NET08_XI829/MM6_d N_XI829/QB_XI829/MM6_g N_VDD_XI829/MM6_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI829/MM5 N_XI829/Q_XI829/MM5_d N_XI829/QB_XI829/MM5_g N_VDD_XI829/MM5_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI829/MM4 N_XI829/QB_XI829/MM4_d N_XI829/Q_XI829/MM4_g N_VDD_XI829/MM4_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI828/MM8 N_XI828/NET08_XI828/MM8_d N_RWL<2>_XI828/MM8_g N_RBL<0>_XI828/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI828/MM7 N_XI828/NET08_XI828/MM7_d N_XI828/QB_XI828/MM7_g N_GND_XI828/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI828/MM10 N_WBL<0>_XI828/MM10_d N_WWLB<2>_XI828/MM10_g N_XI828/Q_XI828/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI828/MM11 N_WBLB<0>_XI828/MM11_d N_WWLB<2>_XI828/MM11_g
+ N_XI828/QB_XI828/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI828/MM1 N_XI828/Q_XI828/MM1_d N_XI828/QB_XI828/MM1_g N_GND_XI828/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI828/MM0 N_XI828/QB_XI828/MM0_d N_XI828/Q_XI828/MM0_g N_GND_XI828/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI828/MM9 N_XI828/NET08_XI828/MM9_d N_RWLB<2>_XI828/MM9_g N_RBL<0>_XI828/MM9_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI828/MM6 N_XI828/NET08_XI828/MM6_d N_XI828/QB_XI828/MM6_g N_VDD_XI828/MM6_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI828/MM5 N_XI828/Q_XI828/MM5_d N_XI828/QB_XI828/MM5_g N_VDD_XI828/MM5_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI828/MM4 N_XI828/QB_XI828/MM4_d N_XI828/Q_XI828/MM4_g N_VDD_XI828/MM4_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI827/MM8 N_XI827/NET08_XI827/MM8_d N_RWL<2>_XI827/MM8_g N_RBL<1>_XI827/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI827/MM7 N_XI827/NET08_XI827/MM7_d N_XI827/QB_XI827/MM7_g N_GND_XI827/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI827/MM10 N_WBL<1>_XI827/MM10_d N_WWLB<2>_XI827/MM10_g N_XI827/Q_XI827/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI827/MM11 N_WBLB<1>_XI827/MM11_d N_WWLB<2>_XI827/MM11_g
+ N_XI827/QB_XI827/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI827/MM1 N_XI827/Q_XI827/MM1_d N_XI827/QB_XI827/MM1_g N_GND_XI827/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI827/MM0 N_XI827/QB_XI827/MM0_d N_XI827/Q_XI827/MM0_g N_GND_XI827/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI827/MM9 N_XI827/NET08_XI827/MM9_d N_RWLB<2>_XI827/MM9_g N_RBL<1>_XI827/MM9_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI827/MM6 N_XI827/NET08_XI827/MM6_d N_XI827/QB_XI827/MM6_g N_VDD_XI827/MM6_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI827/MM5 N_XI827/Q_XI827/MM5_d N_XI827/QB_XI827/MM5_g N_VDD_XI827/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI827/MM4 N_XI827/QB_XI827/MM4_d N_XI827/Q_XI827/MM4_g N_VDD_XI827/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI826/MM8 N_XI826/NET08_XI826/MM8_d N_RWL<2>_XI826/MM8_g N_RBL<2>_XI826/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI826/MM7 N_XI826/NET08_XI826/MM7_d N_XI826/QB_XI826/MM7_g N_GND_XI826/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI826/MM10 N_WBL<2>_XI826/MM10_d N_WWLB<2>_XI826/MM10_g N_XI826/Q_XI826/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI826/MM11 N_WBLB<2>_XI826/MM11_d N_WWLB<2>_XI826/MM11_g
+ N_XI826/QB_XI826/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI826/MM1 N_XI826/Q_XI826/MM1_d N_XI826/QB_XI826/MM1_g N_GND_XI826/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI826/MM0 N_XI826/QB_XI826/MM0_d N_XI826/Q_XI826/MM0_g N_GND_XI826/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI826/MM9 N_XI826/NET08_XI826/MM9_d N_RWLB<2>_XI826/MM9_g N_RBL<2>_XI826/MM9_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI826/MM6 N_XI826/NET08_XI826/MM6_d N_XI826/QB_XI826/MM6_g N_VDD_XI826/MM6_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI826/MM5 N_XI826/Q_XI826/MM5_d N_XI826/QB_XI826/MM5_g N_VDD_XI826/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI826/MM4 N_XI826/QB_XI826/MM4_d N_XI826/Q_XI826/MM4_g N_VDD_XI826/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI850/MM8 N_XI850/NET08_XI850/MM8_d N_RWL<4>_XI850/MM8_g N_RBL<10>_XI850/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI850/MM7 N_XI850/NET08_XI850/MM7_d N_XI850/QB_XI850/MM7_g N_GND_XI850/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI850/MM10 N_WBL<10>_XI850/MM10_d N_WWLB<4>_XI850/MM10_g N_XI850/Q_XI850/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI850/MM11 N_WBLB<10>_XI850/MM11_d N_WWLB<4>_XI850/MM11_g
+ N_XI850/QB_XI850/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI850/MM1 N_XI850/Q_XI850/MM1_d N_XI850/QB_XI850/MM1_g N_GND_XI850/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI850/MM0 N_XI850/QB_XI850/MM0_d N_XI850/Q_XI850/MM0_g N_GND_XI850/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI850/MM9 N_XI850/NET08_XI850/MM9_d N_RWLB<4>_XI850/MM9_g N_RBL<10>_XI850/MM9_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI850/MM6 N_XI850/NET08_XI850/MM6_d N_XI850/QB_XI850/MM6_g N_VDD_XI850/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI850/MM5 N_XI850/Q_XI850/MM5_d N_XI850/QB_XI850/MM5_g N_VDD_XI850/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI850/MM4 N_XI850/QB_XI850/MM4_d N_XI850/Q_XI850/MM4_g N_VDD_XI850/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI849/MM8 N_XI849/NET08_XI849/MM8_d N_RWL<4>_XI849/MM8_g N_RBL<11>_XI849/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI849/MM7 N_XI849/NET08_XI849/MM7_d N_XI849/QB_XI849/MM7_g N_GND_XI849/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI849/MM10 N_WBL<11>_XI849/MM10_d N_WWLB<4>_XI849/MM10_g N_XI849/Q_XI849/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI849/MM11 N_WBLB<11>_XI849/MM11_d N_WWLB<4>_XI849/MM11_g
+ N_XI849/QB_XI849/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI849/MM1 N_XI849/Q_XI849/MM1_d N_XI849/QB_XI849/MM1_g N_GND_XI849/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI849/MM0 N_XI849/QB_XI849/MM0_d N_XI849/Q_XI849/MM0_g N_GND_XI849/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI849/MM9 N_XI849/NET08_XI849/MM9_d N_RWLB<4>_XI849/MM9_g N_RBL<11>_XI849/MM9_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI849/MM6 N_XI849/NET08_XI849/MM6_d N_XI849/QB_XI849/MM6_g N_VDD_XI849/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI849/MM5 N_XI849/Q_XI849/MM5_d N_XI849/QB_XI849/MM5_g N_VDD_XI849/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI849/MM4 N_XI849/QB_XI849/MM4_d N_XI849/Q_XI849/MM4_g N_VDD_XI849/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI848/MM8 N_XI848/NET08_XI848/MM8_d N_RWL<4>_XI848/MM8_g N_RBL<12>_XI848/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI848/MM7 N_XI848/NET08_XI848/MM7_d N_XI848/QB_XI848/MM7_g N_GND_XI848/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI848/MM10 N_WBL<12>_XI848/MM10_d N_WWLB<4>_XI848/MM10_g N_XI848/Q_XI848/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI848/MM11 N_WBLB<12>_XI848/MM11_d N_WWLB<4>_XI848/MM11_g
+ N_XI848/QB_XI848/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI848/MM1 N_XI848/Q_XI848/MM1_d N_XI848/QB_XI848/MM1_g N_GND_XI848/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI848/MM0 N_XI848/QB_XI848/MM0_d N_XI848/Q_XI848/MM0_g N_GND_XI848/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI848/MM9 N_XI848/NET08_XI848/MM9_d N_RWLB<4>_XI848/MM9_g N_RBL<12>_XI848/MM9_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI848/MM6 N_XI848/NET08_XI848/MM6_d N_XI848/QB_XI848/MM6_g N_VDD_XI848/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI848/MM5 N_XI848/Q_XI848/MM5_d N_XI848/QB_XI848/MM5_g N_VDD_XI848/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI848/MM4 N_XI848/QB_XI848/MM4_d N_XI848/Q_XI848/MM4_g N_VDD_XI848/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI851/MM8 N_XI851/NET08_XI851/MM8_d N_RWL<4>_XI851/MM8_g N_RBL<9>_XI851/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI851/MM7 N_XI851/NET08_XI851/MM7_d N_XI851/QB_XI851/MM7_g N_GND_XI851/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI851/MM10 N_WBL<9>_XI851/MM10_d N_WWLB<4>_XI851/MM10_g N_XI851/Q_XI851/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI851/MM11 N_WBLB<9>_XI851/MM11_d N_WWLB<4>_XI851/MM11_g
+ N_XI851/QB_XI851/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI851/MM1 N_XI851/Q_XI851/MM1_d N_XI851/QB_XI851/MM1_g N_GND_XI851/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI851/MM0 N_XI851/QB_XI851/MM0_d N_XI851/Q_XI851/MM0_g N_GND_XI851/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI851/MM9 N_XI851/NET08_XI851/MM9_d N_RWLB<4>_XI851/MM9_g N_RBL<9>_XI851/MM9_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI851/MM6 N_XI851/NET08_XI851/MM6_d N_XI851/QB_XI851/MM6_g N_VDD_XI851/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI851/MM5 N_XI851/Q_XI851/MM5_d N_XI851/QB_XI851/MM5_g N_VDD_XI851/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI851/MM4 N_XI851/QB_XI851/MM4_d N_XI851/Q_XI851/MM4_g N_VDD_XI851/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1026/MM8 N_XI1026/NET08_XI1026/MM8_d N_RWL<15>_XI1026/MM8_g
+ N_RBL<10>_XI1026/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1026/MM7 N_XI1026/NET08_XI1026/MM7_d N_XI1026/QB_XI1026/MM7_g
+ N_GND_XI1026/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1026/MM10 N_WBL<10>_XI1026/MM10_d N_WWLB<15>_XI1026/MM10_g
+ N_XI1026/Q_XI1026/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1026/MM11 N_WBLB<10>_XI1026/MM11_d N_WWLB<15>_XI1026/MM11_g
+ N_XI1026/QB_XI1026/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1026/MM1 N_XI1026/Q_XI1026/MM1_d N_XI1026/QB_XI1026/MM1_g N_GND_XI1026/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1026/MM0 N_XI1026/QB_XI1026/MM0_d N_XI1026/Q_XI1026/MM0_g N_GND_XI1026/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1026/MM9 N_XI1026/NET08_XI1026/MM9_d N_RWLB<15>_XI1026/MM9_g
+ N_RBL<10>_XI1026/MM9_s N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1026/MM6 N_XI1026/NET08_XI1026/MM6_d N_XI1026/QB_XI1026/MM6_g
+ N_VDD_XI1026/MM6_s N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1026/MM5 N_XI1026/Q_XI1026/MM5_d N_XI1026/QB_XI1026/MM5_g N_VDD_XI1026/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1026/MM4 N_XI1026/QB_XI1026/MM4_d N_XI1026/Q_XI1026/MM4_g N_VDD_XI1026/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1001/MM8 N_XI1001/NET08_XI1001/MM8_d N_RWL<13>_XI1001/MM8_g
+ N_RBL<3>_XI1001/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1001/MM7 N_XI1001/NET08_XI1001/MM7_d N_XI1001/QB_XI1001/MM7_g
+ N_GND_XI1001/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1001/MM10 N_WBL<3>_XI1001/MM10_d N_WWLB<13>_XI1001/MM10_g
+ N_XI1001/Q_XI1001/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1001/MM11 N_WBLB<3>_XI1001/MM11_d N_WWLB<13>_XI1001/MM11_g
+ N_XI1001/QB_XI1001/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1001/MM1 N_XI1001/Q_XI1001/MM1_d N_XI1001/QB_XI1001/MM1_g N_GND_XI1001/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1001/MM0 N_XI1001/QB_XI1001/MM0_d N_XI1001/Q_XI1001/MM0_g N_GND_XI1001/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1001/MM9 N_XI1001/NET08_XI1001/MM9_d N_RWLB<13>_XI1001/MM9_g
+ N_RBL<3>_XI1001/MM9_s N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1001/MM6 N_XI1001/NET08_XI1001/MM6_d N_XI1001/QB_XI1001/MM6_g
+ N_VDD_XI1001/MM6_s N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1001/MM5 N_XI1001/Q_XI1001/MM5_d N_XI1001/QB_XI1001/MM5_g N_VDD_XI1001/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1001/MM4 N_XI1001/QB_XI1001/MM4_d N_XI1001/Q_XI1001/MM4_g N_VDD_XI1001/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI854/MM8 N_XI854/NET08_XI854/MM8_d N_RWL<4>_XI854/MM8_g N_RBL<6>_XI854/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI854/MM7 N_XI854/NET08_XI854/MM7_d N_XI854/QB_XI854/MM7_g N_GND_XI854/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI854/MM10 N_WBL<6>_XI854/MM10_d N_WWLB<4>_XI854/MM10_g N_XI854/Q_XI854/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI854/MM11 N_WBLB<6>_XI854/MM11_d N_WWLB<4>_XI854/MM11_g
+ N_XI854/QB_XI854/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI854/MM1 N_XI854/Q_XI854/MM1_d N_XI854/QB_XI854/MM1_g N_GND_XI854/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI854/MM0 N_XI854/QB_XI854/MM0_d N_XI854/Q_XI854/MM0_g N_GND_XI854/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI854/MM9 N_XI854/NET08_XI854/MM9_d N_RWLB<4>_XI854/MM9_g N_RBL<6>_XI854/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI854/MM6 N_XI854/NET08_XI854/MM6_d N_XI854/QB_XI854/MM6_g N_VDD_XI854/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI854/MM5 N_XI854/Q_XI854/MM5_d N_XI854/QB_XI854/MM5_g N_VDD_XI854/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI854/MM4 N_XI854/QB_XI854/MM4_d N_XI854/Q_XI854/MM4_g N_VDD_XI854/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI853/MM8 N_XI853/NET08_XI853/MM8_d N_RWL<4>_XI853/MM8_g N_RBL<7>_XI853/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI853/MM7 N_XI853/NET08_XI853/MM7_d N_XI853/QB_XI853/MM7_g N_GND_XI853/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI853/MM10 N_WBL<7>_XI853/MM10_d N_WWLB<4>_XI853/MM10_g N_XI853/Q_XI853/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI853/MM11 N_WBLB<7>_XI853/MM11_d N_WWLB<4>_XI853/MM11_g
+ N_XI853/QB_XI853/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI853/MM1 N_XI853/Q_XI853/MM1_d N_XI853/QB_XI853/MM1_g N_GND_XI853/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI853/MM0 N_XI853/QB_XI853/MM0_d N_XI853/Q_XI853/MM0_g N_GND_XI853/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI853/MM9 N_XI853/NET08_XI853/MM9_d N_RWLB<4>_XI853/MM9_g N_RBL<7>_XI853/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI853/MM6 N_XI853/NET08_XI853/MM6_d N_XI853/QB_XI853/MM6_g N_VDD_XI853/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI853/MM5 N_XI853/Q_XI853/MM5_d N_XI853/QB_XI853/MM5_g N_VDD_XI853/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI853/MM4 N_XI853/QB_XI853/MM4_d N_XI853/Q_XI853/MM4_g N_VDD_XI853/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI852/MM8 N_XI852/NET08_XI852/MM8_d N_RWL<4>_XI852/MM8_g N_RBL<8>_XI852/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI852/MM7 N_XI852/NET08_XI852/MM7_d N_XI852/QB_XI852/MM7_g N_GND_XI852/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI852/MM10 N_WBL<8>_XI852/MM10_d N_WWLB<4>_XI852/MM10_g N_XI852/Q_XI852/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI852/MM11 N_WBLB<8>_XI852/MM11_d N_WWLB<4>_XI852/MM11_g
+ N_XI852/QB_XI852/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI852/MM1 N_XI852/Q_XI852/MM1_d N_XI852/QB_XI852/MM1_g N_GND_XI852/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI852/MM0 N_XI852/QB_XI852/MM0_d N_XI852/Q_XI852/MM0_g N_GND_XI852/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI852/MM9 N_XI852/NET08_XI852/MM9_d N_RWLB<4>_XI852/MM9_g N_RBL<8>_XI852/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI852/MM6 N_XI852/NET08_XI852/MM6_d N_XI852/QB_XI852/MM6_g N_VDD_XI852/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI852/MM5 N_XI852/Q_XI852/MM5_d N_XI852/QB_XI852/MM5_g N_VDD_XI852/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI852/MM4 N_XI852/QB_XI852/MM4_d N_XI852/Q_XI852/MM4_g N_VDD_XI852/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI855/MM8 N_XI855/NET08_XI855/MM8_d N_RWL<4>_XI855/MM8_g N_RBL<5>_XI855/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI855/MM7 N_XI855/NET08_XI855/MM7_d N_XI855/QB_XI855/MM7_g N_GND_XI855/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI855/MM10 N_WBL<5>_XI855/MM10_d N_WWLB<4>_XI855/MM10_g N_XI855/Q_XI855/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI855/MM11 N_WBLB<5>_XI855/MM11_d N_WWLB<4>_XI855/MM11_g
+ N_XI855/QB_XI855/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI855/MM1 N_XI855/Q_XI855/MM1_d N_XI855/QB_XI855/MM1_g N_GND_XI855/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI855/MM0 N_XI855/QB_XI855/MM0_d N_XI855/Q_XI855/MM0_g N_GND_XI855/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI855/MM9 N_XI855/NET08_XI855/MM9_d N_RWLB<4>_XI855/MM9_g N_RBL<5>_XI855/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI855/MM6 N_XI855/NET08_XI855/MM6_d N_XI855/QB_XI855/MM6_g N_VDD_XI855/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI855/MM5 N_XI855/Q_XI855/MM5_d N_XI855/QB_XI855/MM5_g N_VDD_XI855/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI855/MM4 N_XI855/QB_XI855/MM4_d N_XI855/Q_XI855/MM4_g N_VDD_XI855/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI880/MM8 N_XI880/NET08_XI880/MM8_d N_RWL<6>_XI880/MM8_g N_RBL<12>_XI880/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI880/MM7 N_XI880/NET08_XI880/MM7_d N_XI880/QB_XI880/MM7_g N_GND_XI880/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI880/MM10 N_WBL<12>_XI880/MM10_d N_WWLB<6>_XI880/MM10_g N_XI880/Q_XI880/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI880/MM11 N_WBLB<12>_XI880/MM11_d N_WWLB<6>_XI880/MM11_g
+ N_XI880/QB_XI880/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI880/MM1 N_XI880/Q_XI880/MM1_d N_XI880/QB_XI880/MM1_g N_GND_XI880/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI880/MM0 N_XI880/QB_XI880/MM0_d N_XI880/Q_XI880/MM0_g N_GND_XI880/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI880/MM9 N_XI880/NET08_XI880/MM9_d N_RWLB<6>_XI880/MM9_g N_RBL<12>_XI880/MM9_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI880/MM6 N_XI880/NET08_XI880/MM6_d N_XI880/QB_XI880/MM6_g N_VDD_XI880/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI880/MM5 N_XI880/Q_XI880/MM5_d N_XI880/QB_XI880/MM5_g N_VDD_XI880/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI880/MM4 N_XI880/QB_XI880/MM4_d N_XI880/Q_XI880/MM4_g N_VDD_XI880/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI794/MM8 N_XI794/NET08_XI794/MM8_d N_RWL<0>_XI794/MM8_g N_RBL<3>_XI794/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI794/MM7 N_XI794/NET08_XI794/MM7_d N_XI794/QB_XI794/MM7_g N_GND_XI794/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI794/MM10 N_WBL<3>_XI794/MM10_d N_WWLB<0>_XI794/MM10_g N_XI794/Q_XI794/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI794/MM11 N_WBLB<3>_XI794/MM11_d N_WWLB<0>_XI794/MM11_g
+ N_XI794/QB_XI794/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI794/MM1 N_XI794/Q_XI794/MM1_d N_XI794/QB_XI794/MM1_g N_GND_XI794/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI794/MM0 N_XI794/QB_XI794/MM0_d N_XI794/Q_XI794/MM0_g N_GND_XI794/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI794/MM9 N_XI794/NET08_XI794/MM9_d N_RWLB<0>_XI794/MM9_g N_RBL<3>_XI794/MM9_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI794/MM6 N_XI794/NET08_XI794/MM6_d N_XI794/QB_XI794/MM6_g N_VDD_XI794/MM6_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI794/MM5 N_XI794/Q_XI794/MM5_d N_XI794/QB_XI794/MM5_g N_VDD_XI794/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI794/MM4 N_XI794/QB_XI794/MM4_d N_XI794/Q_XI794/MM4_g N_VDD_XI794/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI825/MM8 N_XI825/NET08_XI825/MM8_d N_RWL<2>_XI825/MM8_g N_RBL<3>_XI825/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI825/MM7 N_XI825/NET08_XI825/MM7_d N_XI825/QB_XI825/MM7_g N_GND_XI825/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI825/MM10 N_WBL<3>_XI825/MM10_d N_WWLB<2>_XI825/MM10_g N_XI825/Q_XI825/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI825/MM11 N_WBLB<3>_XI825/MM11_d N_WWLB<2>_XI825/MM11_g
+ N_XI825/QB_XI825/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI825/MM1 N_XI825/Q_XI825/MM1_d N_XI825/QB_XI825/MM1_g N_GND_XI825/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI825/MM0 N_XI825/QB_XI825/MM0_d N_XI825/Q_XI825/MM0_g N_GND_XI825/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI825/MM9 N_XI825/NET08_XI825/MM9_d N_RWLB<2>_XI825/MM9_g N_RBL<3>_XI825/MM9_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI825/MM6 N_XI825/NET08_XI825/MM6_d N_XI825/QB_XI825/MM6_g N_VDD_XI825/MM6_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI825/MM5 N_XI825/Q_XI825/MM5_d N_XI825/QB_XI825/MM5_g N_VDD_XI825/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI825/MM4 N_XI825/QB_XI825/MM4_d N_XI825/Q_XI825/MM4_g N_VDD_XI825/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI824/MM8 N_XI824/NET08_XI824/MM8_d N_RWL<2>_XI824/MM8_g N_RBL<4>_XI824/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI824/MM7 N_XI824/NET08_XI824/MM7_d N_XI824/QB_XI824/MM7_g N_GND_XI824/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI824/MM10 N_WBL<4>_XI824/MM10_d N_WWLB<2>_XI824/MM10_g N_XI824/Q_XI824/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI824/MM11 N_WBLB<4>_XI824/MM11_d N_WWLB<2>_XI824/MM11_g
+ N_XI824/QB_XI824/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI824/MM1 N_XI824/Q_XI824/MM1_d N_XI824/QB_XI824/MM1_g N_GND_XI824/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI824/MM0 N_XI824/QB_XI824/MM0_d N_XI824/Q_XI824/MM0_g N_GND_XI824/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI824/MM9 N_XI824/NET08_XI824/MM9_d N_RWLB<2>_XI824/MM9_g N_RBL<4>_XI824/MM9_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI824/MM6 N_XI824/NET08_XI824/MM6_d N_XI824/QB_XI824/MM6_g N_VDD_XI824/MM6_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI824/MM5 N_XI824/Q_XI824/MM5_d N_XI824/QB_XI824/MM5_g N_VDD_XI824/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI824/MM4 N_XI824/QB_XI824/MM4_d N_XI824/Q_XI824/MM4_g N_VDD_XI824/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI823/MM8 N_XI823/NET08_XI823/MM8_d N_RWL<2>_XI823/MM8_g N_RBL<5>_XI823/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI823/MM7 N_XI823/NET08_XI823/MM7_d N_XI823/QB_XI823/MM7_g N_GND_XI823/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI823/MM10 N_WBL<5>_XI823/MM10_d N_WWLB<2>_XI823/MM10_g N_XI823/Q_XI823/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI823/MM11 N_WBLB<5>_XI823/MM11_d N_WWLB<2>_XI823/MM11_g
+ N_XI823/QB_XI823/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI823/MM1 N_XI823/Q_XI823/MM1_d N_XI823/QB_XI823/MM1_g N_GND_XI823/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI823/MM0 N_XI823/QB_XI823/MM0_d N_XI823/Q_XI823/MM0_g N_GND_XI823/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI823/MM9 N_XI823/NET08_XI823/MM9_d N_RWLB<2>_XI823/MM9_g N_RBL<5>_XI823/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI823/MM6 N_XI823/NET08_XI823/MM6_d N_XI823/QB_XI823/MM6_g N_VDD_XI823/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI823/MM5 N_XI823/Q_XI823/MM5_d N_XI823/QB_XI823/MM5_g N_VDD_XI823/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI823/MM4 N_XI823/QB_XI823/MM4_d N_XI823/Q_XI823/MM4_g N_VDD_XI823/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI822/MM8 N_XI822/NET08_XI822/MM8_d N_RWL<2>_XI822/MM8_g N_RBL<6>_XI822/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI822/MM7 N_XI822/NET08_XI822/MM7_d N_XI822/QB_XI822/MM7_g N_GND_XI822/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI822/MM10 N_WBL<6>_XI822/MM10_d N_WWLB<2>_XI822/MM10_g N_XI822/Q_XI822/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI822/MM11 N_WBLB<6>_XI822/MM11_d N_WWLB<2>_XI822/MM11_g
+ N_XI822/QB_XI822/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI822/MM1 N_XI822/Q_XI822/MM1_d N_XI822/QB_XI822/MM1_g N_GND_XI822/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI822/MM0 N_XI822/QB_XI822/MM0_d N_XI822/Q_XI822/MM0_g N_GND_XI822/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI822/MM9 N_XI822/NET08_XI822/MM9_d N_RWLB<2>_XI822/MM9_g N_RBL<6>_XI822/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI822/MM6 N_XI822/NET08_XI822/MM6_d N_XI822/QB_XI822/MM6_g N_VDD_XI822/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI822/MM5 N_XI822/Q_XI822/MM5_d N_XI822/QB_XI822/MM5_g N_VDD_XI822/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI822/MM4 N_XI822/QB_XI822/MM4_d N_XI822/Q_XI822/MM4_g N_VDD_XI822/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI821/MM8 N_XI821/NET08_XI821/MM8_d N_RWL<2>_XI821/MM8_g N_RBL<7>_XI821/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI821/MM7 N_XI821/NET08_XI821/MM7_d N_XI821/QB_XI821/MM7_g N_GND_XI821/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI821/MM10 N_WBL<7>_XI821/MM10_d N_WWLB<2>_XI821/MM10_g N_XI821/Q_XI821/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI821/MM11 N_WBLB<7>_XI821/MM11_d N_WWLB<2>_XI821/MM11_g
+ N_XI821/QB_XI821/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI821/MM1 N_XI821/Q_XI821/MM1_d N_XI821/QB_XI821/MM1_g N_GND_XI821/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI821/MM0 N_XI821/QB_XI821/MM0_d N_XI821/Q_XI821/MM0_g N_GND_XI821/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI821/MM9 N_XI821/NET08_XI821/MM9_d N_RWLB<2>_XI821/MM9_g N_RBL<7>_XI821/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI821/MM6 N_XI821/NET08_XI821/MM6_d N_XI821/QB_XI821/MM6_g N_VDD_XI821/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI821/MM5 N_XI821/Q_XI821/MM5_d N_XI821/QB_XI821/MM5_g N_VDD_XI821/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI821/MM4 N_XI821/QB_XI821/MM4_d N_XI821/Q_XI821/MM4_g N_VDD_XI821/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI820/MM8 N_XI820/NET08_XI820/MM8_d N_RWL<2>_XI820/MM8_g N_RBL<8>_XI820/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI820/MM7 N_XI820/NET08_XI820/MM7_d N_XI820/QB_XI820/MM7_g N_GND_XI820/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI820/MM10 N_WBL<8>_XI820/MM10_d N_WWLB<2>_XI820/MM10_g N_XI820/Q_XI820/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI820/MM11 N_WBLB<8>_XI820/MM11_d N_WWLB<2>_XI820/MM11_g
+ N_XI820/QB_XI820/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI820/MM1 N_XI820/Q_XI820/MM1_d N_XI820/QB_XI820/MM1_g N_GND_XI820/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI820/MM0 N_XI820/QB_XI820/MM0_d N_XI820/Q_XI820/MM0_g N_GND_XI820/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI820/MM9 N_XI820/NET08_XI820/MM9_d N_RWLB<2>_XI820/MM9_g N_RBL<8>_XI820/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI820/MM6 N_XI820/NET08_XI820/MM6_d N_XI820/QB_XI820/MM6_g N_VDD_XI820/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI820/MM5 N_XI820/Q_XI820/MM5_d N_XI820/QB_XI820/MM5_g N_VDD_XI820/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI820/MM4 N_XI820/QB_XI820/MM4_d N_XI820/Q_XI820/MM4_g N_VDD_XI820/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI847/MM8 N_XI847/NET08_XI847/MM8_d N_RWL<4>_XI847/MM8_g N_RBL<13>_XI847/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI847/MM7 N_XI847/NET08_XI847/MM7_d N_XI847/QB_XI847/MM7_g N_GND_XI847/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI847/MM10 N_WBL<13>_XI847/MM10_d N_WWLB<4>_XI847/MM10_g N_XI847/Q_XI847/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI847/MM11 N_WBLB<13>_XI847/MM11_d N_WWLB<4>_XI847/MM11_g
+ N_XI847/QB_XI847/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI847/MM1 N_XI847/Q_XI847/MM1_d N_XI847/QB_XI847/MM1_g N_GND_XI847/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI847/MM0 N_XI847/QB_XI847/MM0_d N_XI847/Q_XI847/MM0_g N_GND_XI847/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI847/MM9 N_XI847/NET08_XI847/MM9_d N_RWLB<4>_XI847/MM9_g N_RBL<13>_XI847/MM9_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI847/MM6 N_XI847/NET08_XI847/MM6_d N_XI847/QB_XI847/MM6_g N_VDD_XI847/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI847/MM5 N_XI847/Q_XI847/MM5_d N_XI847/QB_XI847/MM5_g N_VDD_XI847/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI847/MM4 N_XI847/QB_XI847/MM4_d N_XI847/Q_XI847/MM4_g N_VDD_XI847/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI846/MM8 N_XI846/NET08_XI846/MM8_d N_RWL<4>_XI846/MM8_g N_RBL<14>_XI846/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI846/MM7 N_XI846/NET08_XI846/MM7_d N_XI846/QB_XI846/MM7_g N_GND_XI846/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI846/MM10 N_WBL<14>_XI846/MM10_d N_WWLB<4>_XI846/MM10_g N_XI846/Q_XI846/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI846/MM11 N_WBLB<14>_XI846/MM11_d N_WWLB<4>_XI846/MM11_g
+ N_XI846/QB_XI846/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI846/MM1 N_XI846/Q_XI846/MM1_d N_XI846/QB_XI846/MM1_g N_GND_XI846/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI846/MM0 N_XI846/QB_XI846/MM0_d N_XI846/Q_XI846/MM0_g N_GND_XI846/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI846/MM9 N_XI846/NET08_XI846/MM9_d N_RWLB<4>_XI846/MM9_g N_RBL<14>_XI846/MM9_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI846/MM6 N_XI846/NET08_XI846/MM6_d N_XI846/QB_XI846/MM6_g N_VDD_XI846/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI846/MM5 N_XI846/Q_XI846/MM5_d N_XI846/QB_XI846/MM5_g N_VDD_XI846/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI846/MM4 N_XI846/QB_XI846/MM4_d N_XI846/Q_XI846/MM4_g N_VDD_XI846/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI845/MM8 N_XI845/NET08_XI845/MM8_d N_RWL<3>_XI845/MM8_g N_RBL<15>_XI845/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI845/MM7 N_XI845/NET08_XI845/MM7_d N_XI845/QB_XI845/MM7_g N_GND_XI845/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI845/MM10 N_WBL<15>_XI845/MM10_d N_WWLB<3>_XI845/MM10_g N_XI845/Q_XI845/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI845/MM11 N_WBLB<15>_XI845/MM11_d N_WWLB<3>_XI845/MM11_g
+ N_XI845/QB_XI845/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI845/MM1 N_XI845/Q_XI845/MM1_d N_XI845/QB_XI845/MM1_g N_GND_XI845/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI845/MM0 N_XI845/QB_XI845/MM0_d N_XI845/Q_XI845/MM0_g N_GND_XI845/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI845/MM9 N_XI845/NET08_XI845/MM9_d N_RWLB<3>_XI845/MM9_g N_RBL<15>_XI845/MM9_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI845/MM6 N_XI845/NET08_XI845/MM6_d N_XI845/QB_XI845/MM6_g N_VDD_XI845/MM6_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI845/MM5 N_XI845/Q_XI845/MM5_d N_XI845/QB_XI845/MM5_g N_VDD_XI845/MM5_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI845/MM4 N_XI845/QB_XI845/MM4_d N_XI845/Q_XI845/MM4_g N_VDD_XI845/MM4_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI844/MM8 N_XI844/NET08_XI844/MM8_d N_RWL<3>_XI844/MM8_g N_RBL<0>_XI844/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI844/MM7 N_XI844/NET08_XI844/MM7_d N_XI844/QB_XI844/MM7_g N_GND_XI844/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI844/MM10 N_WBL<0>_XI844/MM10_d N_WWLB<3>_XI844/MM10_g N_XI844/Q_XI844/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI844/MM11 N_WBLB<0>_XI844/MM11_d N_WWLB<3>_XI844/MM11_g
+ N_XI844/QB_XI844/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI844/MM1 N_XI844/Q_XI844/MM1_d N_XI844/QB_XI844/MM1_g N_GND_XI844/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI844/MM0 N_XI844/QB_XI844/MM0_d N_XI844/Q_XI844/MM0_g N_GND_XI844/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI844/MM9 N_XI844/NET08_XI844/MM9_d N_RWLB<3>_XI844/MM9_g N_RBL<0>_XI844/MM9_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI844/MM6 N_XI844/NET08_XI844/MM6_d N_XI844/QB_XI844/MM6_g N_VDD_XI844/MM6_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI844/MM5 N_XI844/Q_XI844/MM5_d N_XI844/QB_XI844/MM5_g N_VDD_XI844/MM5_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI844/MM4 N_XI844/QB_XI844/MM4_d N_XI844/Q_XI844/MM4_g N_VDD_XI844/MM4_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1025/MM8 N_XI1025/NET08_XI1025/MM8_d N_RWL<15>_XI1025/MM8_g
+ N_RBL<11>_XI1025/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1025/MM7 N_XI1025/NET08_XI1025/MM7_d N_XI1025/QB_XI1025/MM7_g
+ N_GND_XI1025/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1025/MM10 N_WBL<11>_XI1025/MM10_d N_WWLB<15>_XI1025/MM10_g
+ N_XI1025/Q_XI1025/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1025/MM11 N_WBLB<11>_XI1025/MM11_d N_WWLB<15>_XI1025/MM11_g
+ N_XI1025/QB_XI1025/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1025/MM1 N_XI1025/Q_XI1025/MM1_d N_XI1025/QB_XI1025/MM1_g N_GND_XI1025/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1025/MM0 N_XI1025/QB_XI1025/MM0_d N_XI1025/Q_XI1025/MM0_g N_GND_XI1025/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1025/MM9 N_XI1025/NET08_XI1025/MM9_d N_RWLB<15>_XI1025/MM9_g
+ N_RBL<11>_XI1025/MM9_s N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1025/MM6 N_XI1025/NET08_XI1025/MM6_d N_XI1025/QB_XI1025/MM6_g
+ N_VDD_XI1025/MM6_s N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1025/MM5 N_XI1025/Q_XI1025/MM5_d N_XI1025/QB_XI1025/MM5_g N_VDD_XI1025/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1025/MM4 N_XI1025/QB_XI1025/MM4_d N_XI1025/Q_XI1025/MM4_g N_VDD_XI1025/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1002/MM8 N_XI1002/NET08_XI1002/MM8_d N_RWL<13>_XI1002/MM8_g
+ N_RBL<2>_XI1002/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1002/MM7 N_XI1002/NET08_XI1002/MM7_d N_XI1002/QB_XI1002/MM7_g
+ N_GND_XI1002/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1002/MM10 N_WBL<2>_XI1002/MM10_d N_WWLB<13>_XI1002/MM10_g
+ N_XI1002/Q_XI1002/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1002/MM11 N_WBLB<2>_XI1002/MM11_d N_WWLB<13>_XI1002/MM11_g
+ N_XI1002/QB_XI1002/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1002/MM1 N_XI1002/Q_XI1002/MM1_d N_XI1002/QB_XI1002/MM1_g N_GND_XI1002/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1002/MM0 N_XI1002/QB_XI1002/MM0_d N_XI1002/Q_XI1002/MM0_g N_GND_XI1002/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1002/MM9 N_XI1002/NET08_XI1002/MM9_d N_RWLB<13>_XI1002/MM9_g
+ N_RBL<2>_XI1002/MM9_s N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1002/MM6 N_XI1002/NET08_XI1002/MM6_d N_XI1002/QB_XI1002/MM6_g
+ N_VDD_XI1002/MM6_s N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1002/MM5 N_XI1002/Q_XI1002/MM5_d N_XI1002/QB_XI1002/MM5_g N_VDD_XI1002/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1002/MM4 N_XI1002/QB_XI1002/MM4_d N_XI1002/Q_XI1002/MM4_g N_VDD_XI1002/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI801/MM8 N_XI801/NET08_XI801/MM8_d N_RWL<1>_XI801/MM8_g N_RBL<11>_XI801/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI801/MM7 N_XI801/NET08_XI801/MM7_d N_XI801/QB_XI801/MM7_g N_GND_XI801/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI801/MM10 N_WBL<11>_XI801/MM10_d N_WWLB<1>_XI801/MM10_g N_XI801/Q_XI801/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI801/MM11 N_WBLB<11>_XI801/MM11_d N_WWLB<1>_XI801/MM11_g
+ N_XI801/QB_XI801/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI801/MM1 N_XI801/Q_XI801/MM1_d N_XI801/QB_XI801/MM1_g N_GND_XI801/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI801/MM0 N_XI801/QB_XI801/MM0_d N_XI801/Q_XI801/MM0_g N_GND_XI801/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI801/MM9 N_XI801/NET08_XI801/MM9_d N_RWLB<1>_XI801/MM9_g N_RBL<11>_XI801/MM9_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI801/MM6 N_XI801/NET08_XI801/MM6_d N_XI801/QB_XI801/MM6_g N_VDD_XI801/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI801/MM5 N_XI801/Q_XI801/MM5_d N_XI801/QB_XI801/MM5_g N_VDD_XI801/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI801/MM4 N_XI801/QB_XI801/MM4_d N_XI801/Q_XI801/MM4_g N_VDD_XI801/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI800/MM8 N_XI800/NET08_XI800/MM8_d N_RWL<1>_XI800/MM8_g N_RBL<12>_XI800/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI800/MM7 N_XI800/NET08_XI800/MM7_d N_XI800/QB_XI800/MM7_g N_GND_XI800/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI800/MM10 N_WBL<12>_XI800/MM10_d N_WWLB<1>_XI800/MM10_g N_XI800/Q_XI800/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI800/MM11 N_WBLB<12>_XI800/MM11_d N_WWLB<1>_XI800/MM11_g
+ N_XI800/QB_XI800/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI800/MM1 N_XI800/Q_XI800/MM1_d N_XI800/QB_XI800/MM1_g N_GND_XI800/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI800/MM0 N_XI800/QB_XI800/MM0_d N_XI800/Q_XI800/MM0_g N_GND_XI800/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI800/MM9 N_XI800/NET08_XI800/MM9_d N_RWLB<1>_XI800/MM9_g N_RBL<12>_XI800/MM9_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI800/MM6 N_XI800/NET08_XI800/MM6_d N_XI800/QB_XI800/MM6_g N_VDD_XI800/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI800/MM5 N_XI800/Q_XI800/MM5_d N_XI800/QB_XI800/MM5_g N_VDD_XI800/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI800/MM4 N_XI800/QB_XI800/MM4_d N_XI800/Q_XI800/MM4_g N_VDD_XI800/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI799/MM8 N_XI799/NET08_XI799/MM8_d N_RWL<1>_XI799/MM8_g N_RBL<13>_XI799/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI799/MM7 N_XI799/NET08_XI799/MM7_d N_XI799/QB_XI799/MM7_g N_GND_XI799/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI799/MM10 N_WBL<13>_XI799/MM10_d N_WWLB<1>_XI799/MM10_g N_XI799/Q_XI799/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI799/MM11 N_WBLB<13>_XI799/MM11_d N_WWLB<1>_XI799/MM11_g
+ N_XI799/QB_XI799/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI799/MM1 N_XI799/Q_XI799/MM1_d N_XI799/QB_XI799/MM1_g N_GND_XI799/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI799/MM0 N_XI799/QB_XI799/MM0_d N_XI799/Q_XI799/MM0_g N_GND_XI799/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI799/MM9 N_XI799/NET08_XI799/MM9_d N_RWLB<1>_XI799/MM9_g N_RBL<13>_XI799/MM9_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI799/MM6 N_XI799/NET08_XI799/MM6_d N_XI799/QB_XI799/MM6_g N_VDD_XI799/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI799/MM5 N_XI799/Q_XI799/MM5_d N_XI799/QB_XI799/MM5_g N_VDD_XI799/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI799/MM4 N_XI799/QB_XI799/MM4_d N_XI799/Q_XI799/MM4_g N_VDD_XI799/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI798/MM8 N_XI798/NET08_XI798/MM8_d N_RWL<1>_XI798/MM8_g N_RBL<14>_XI798/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI798/MM7 N_XI798/NET08_XI798/MM7_d N_XI798/QB_XI798/MM7_g N_GND_XI798/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI798/MM10 N_WBL<14>_XI798/MM10_d N_WWLB<1>_XI798/MM10_g N_XI798/Q_XI798/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI798/MM11 N_WBLB<14>_XI798/MM11_d N_WWLB<1>_XI798/MM11_g
+ N_XI798/QB_XI798/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI798/MM1 N_XI798/Q_XI798/MM1_d N_XI798/QB_XI798/MM1_g N_GND_XI798/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI798/MM0 N_XI798/QB_XI798/MM0_d N_XI798/Q_XI798/MM0_g N_GND_XI798/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI798/MM9 N_XI798/NET08_XI798/MM9_d N_RWLB<1>_XI798/MM9_g N_RBL<14>_XI798/MM9_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI798/MM6 N_XI798/NET08_XI798/MM6_d N_XI798/QB_XI798/MM6_g N_VDD_XI798/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI798/MM5 N_XI798/Q_XI798/MM5_d N_XI798/QB_XI798/MM5_g N_VDD_XI798/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI798/MM4 N_XI798/QB_XI798/MM4_d N_XI798/Q_XI798/MM4_g N_VDD_XI798/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI791/MM8 N_XI791/NET08_XI791/MM8_d N_RWL<0>_XI791/MM8_g N_RBL<6>_XI791/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI791/MM7 N_XI791/NET08_XI791/MM7_d N_XI791/QB_XI791/MM7_g N_GND_XI791/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI791/MM10 N_WBL<6>_XI791/MM10_d N_WWLB<0>_XI791/MM10_g N_XI791/Q_XI791/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI791/MM11 N_WBLB<6>_XI791/MM11_d N_WWLB<0>_XI791/MM11_g
+ N_XI791/QB_XI791/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI791/MM1 N_XI791/Q_XI791/MM1_d N_XI791/QB_XI791/MM1_g N_GND_XI791/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI791/MM0 N_XI791/QB_XI791/MM0_d N_XI791/Q_XI791/MM0_g N_GND_XI791/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI791/MM9 N_XI791/NET08_XI791/MM9_d N_RWLB<0>_XI791/MM9_g N_RBL<6>_XI791/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI791/MM6 N_XI791/NET08_XI791/MM6_d N_XI791/QB_XI791/MM6_g N_VDD_XI791/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI791/MM5 N_XI791/Q_XI791/MM5_d N_XI791/QB_XI791/MM5_g N_VDD_XI791/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI791/MM4 N_XI791/QB_XI791/MM4_d N_XI791/Q_XI791/MM4_g N_VDD_XI791/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI790/MM8 N_XI790/NET08_XI790/MM8_d N_RWL<0>_XI790/MM8_g N_RBL<7>_XI790/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI790/MM7 N_XI790/NET08_XI790/MM7_d N_XI790/QB_XI790/MM7_g N_GND_XI790/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI790/MM10 N_WBL<7>_XI790/MM10_d N_WWLB<0>_XI790/MM10_g N_XI790/Q_XI790/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI790/MM11 N_WBLB<7>_XI790/MM11_d N_WWLB<0>_XI790/MM11_g
+ N_XI790/QB_XI790/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI790/MM1 N_XI790/Q_XI790/MM1_d N_XI790/QB_XI790/MM1_g N_GND_XI790/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI790/MM0 N_XI790/QB_XI790/MM0_d N_XI790/Q_XI790/MM0_g N_GND_XI790/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI790/MM9 N_XI790/NET08_XI790/MM9_d N_RWLB<0>_XI790/MM9_g N_RBL<7>_XI790/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI790/MM6 N_XI790/NET08_XI790/MM6_d N_XI790/QB_XI790/MM6_g N_VDD_XI790/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI790/MM5 N_XI790/Q_XI790/MM5_d N_XI790/QB_XI790/MM5_g N_VDD_XI790/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI790/MM4 N_XI790/QB_XI790/MM4_d N_XI790/Q_XI790/MM4_g N_VDD_XI790/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI819/MM8 N_XI819/NET08_XI819/MM8_d N_RWL<2>_XI819/MM8_g N_RBL<9>_XI819/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI819/MM7 N_XI819/NET08_XI819/MM7_d N_XI819/QB_XI819/MM7_g N_GND_XI819/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI819/MM10 N_WBL<9>_XI819/MM10_d N_WWLB<2>_XI819/MM10_g N_XI819/Q_XI819/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI819/MM11 N_WBLB<9>_XI819/MM11_d N_WWLB<2>_XI819/MM11_g
+ N_XI819/QB_XI819/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI819/MM1 N_XI819/Q_XI819/MM1_d N_XI819/QB_XI819/MM1_g N_GND_XI819/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI819/MM0 N_XI819/QB_XI819/MM0_d N_XI819/Q_XI819/MM0_g N_GND_XI819/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI819/MM9 N_XI819/NET08_XI819/MM9_d N_RWLB<2>_XI819/MM9_g N_RBL<9>_XI819/MM9_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI819/MM6 N_XI819/NET08_XI819/MM6_d N_XI819/QB_XI819/MM6_g N_VDD_XI819/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI819/MM5 N_XI819/Q_XI819/MM5_d N_XI819/QB_XI819/MM5_g N_VDD_XI819/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI819/MM4 N_XI819/QB_XI819/MM4_d N_XI819/Q_XI819/MM4_g N_VDD_XI819/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI818/MM8 N_XI818/NET08_XI818/MM8_d N_RWL<2>_XI818/MM8_g N_RBL<10>_XI818/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI818/MM7 N_XI818/NET08_XI818/MM7_d N_XI818/QB_XI818/MM7_g N_GND_XI818/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI818/MM10 N_WBL<10>_XI818/MM10_d N_WWLB<2>_XI818/MM10_g N_XI818/Q_XI818/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI818/MM11 N_WBLB<10>_XI818/MM11_d N_WWLB<2>_XI818/MM11_g
+ N_XI818/QB_XI818/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI818/MM1 N_XI818/Q_XI818/MM1_d N_XI818/QB_XI818/MM1_g N_GND_XI818/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI818/MM0 N_XI818/QB_XI818/MM0_d N_XI818/Q_XI818/MM0_g N_GND_XI818/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI818/MM9 N_XI818/NET08_XI818/MM9_d N_RWLB<2>_XI818/MM9_g N_RBL<10>_XI818/MM9_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI818/MM6 N_XI818/NET08_XI818/MM6_d N_XI818/QB_XI818/MM6_g N_VDD_XI818/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI818/MM5 N_XI818/Q_XI818/MM5_d N_XI818/QB_XI818/MM5_g N_VDD_XI818/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI818/MM4 N_XI818/QB_XI818/MM4_d N_XI818/Q_XI818/MM4_g N_VDD_XI818/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI817/MM8 N_XI817/NET08_XI817/MM8_d N_RWL<2>_XI817/MM8_g N_RBL<11>_XI817/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI817/MM7 N_XI817/NET08_XI817/MM7_d N_XI817/QB_XI817/MM7_g N_GND_XI817/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI817/MM10 N_WBL<11>_XI817/MM10_d N_WWLB<2>_XI817/MM10_g N_XI817/Q_XI817/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI817/MM11 N_WBLB<11>_XI817/MM11_d N_WWLB<2>_XI817/MM11_g
+ N_XI817/QB_XI817/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI817/MM1 N_XI817/Q_XI817/MM1_d N_XI817/QB_XI817/MM1_g N_GND_XI817/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI817/MM0 N_XI817/QB_XI817/MM0_d N_XI817/Q_XI817/MM0_g N_GND_XI817/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI817/MM9 N_XI817/NET08_XI817/MM9_d N_RWLB<2>_XI817/MM9_g N_RBL<11>_XI817/MM9_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI817/MM6 N_XI817/NET08_XI817/MM6_d N_XI817/QB_XI817/MM6_g N_VDD_XI817/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI817/MM5 N_XI817/Q_XI817/MM5_d N_XI817/QB_XI817/MM5_g N_VDD_XI817/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI817/MM4 N_XI817/QB_XI817/MM4_d N_XI817/Q_XI817/MM4_g N_VDD_XI817/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI816/MM8 N_XI816/NET08_XI816/MM8_d N_RWL<2>_XI816/MM8_g N_RBL<12>_XI816/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI816/MM7 N_XI816/NET08_XI816/MM7_d N_XI816/QB_XI816/MM7_g N_GND_XI816/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI816/MM10 N_WBL<12>_XI816/MM10_d N_WWLB<2>_XI816/MM10_g N_XI816/Q_XI816/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI816/MM11 N_WBLB<12>_XI816/MM11_d N_WWLB<2>_XI816/MM11_g
+ N_XI816/QB_XI816/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI816/MM1 N_XI816/Q_XI816/MM1_d N_XI816/QB_XI816/MM1_g N_GND_XI816/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI816/MM0 N_XI816/QB_XI816/MM0_d N_XI816/Q_XI816/MM0_g N_GND_XI816/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI816/MM9 N_XI816/NET08_XI816/MM9_d N_RWLB<2>_XI816/MM9_g N_RBL<12>_XI816/MM9_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI816/MM6 N_XI816/NET08_XI816/MM6_d N_XI816/QB_XI816/MM6_g N_VDD_XI816/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI816/MM5 N_XI816/Q_XI816/MM5_d N_XI816/QB_XI816/MM5_g N_VDD_XI816/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI816/MM4 N_XI816/QB_XI816/MM4_d N_XI816/Q_XI816/MM4_g N_VDD_XI816/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI815/MM8 N_XI815/NET08_XI815/MM8_d N_RWL<2>_XI815/MM8_g N_RBL<13>_XI815/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI815/MM7 N_XI815/NET08_XI815/MM7_d N_XI815/QB_XI815/MM7_g N_GND_XI815/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI815/MM10 N_WBL<13>_XI815/MM10_d N_WWLB<2>_XI815/MM10_g N_XI815/Q_XI815/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI815/MM11 N_WBLB<13>_XI815/MM11_d N_WWLB<2>_XI815/MM11_g
+ N_XI815/QB_XI815/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI815/MM1 N_XI815/Q_XI815/MM1_d N_XI815/QB_XI815/MM1_g N_GND_XI815/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI815/MM0 N_XI815/QB_XI815/MM0_d N_XI815/Q_XI815/MM0_g N_GND_XI815/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI815/MM9 N_XI815/NET08_XI815/MM9_d N_RWLB<2>_XI815/MM9_g N_RBL<13>_XI815/MM9_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI815/MM6 N_XI815/NET08_XI815/MM6_d N_XI815/QB_XI815/MM6_g N_VDD_XI815/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI815/MM5 N_XI815/Q_XI815/MM5_d N_XI815/QB_XI815/MM5_g N_VDD_XI815/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI815/MM4 N_XI815/QB_XI815/MM4_d N_XI815/Q_XI815/MM4_g N_VDD_XI815/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI814/MM8 N_XI814/NET08_XI814/MM8_d N_RWL<2>_XI814/MM8_g N_RBL<14>_XI814/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI814/MM7 N_XI814/NET08_XI814/MM7_d N_XI814/QB_XI814/MM7_g N_GND_XI814/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI814/MM10 N_WBL<14>_XI814/MM10_d N_WWLB<2>_XI814/MM10_g N_XI814/Q_XI814/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI814/MM11 N_WBLB<14>_XI814/MM11_d N_WWLB<2>_XI814/MM11_g
+ N_XI814/QB_XI814/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI814/MM1 N_XI814/Q_XI814/MM1_d N_XI814/QB_XI814/MM1_g N_GND_XI814/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI814/MM0 N_XI814/QB_XI814/MM0_d N_XI814/Q_XI814/MM0_g N_GND_XI814/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI814/MM9 N_XI814/NET08_XI814/MM9_d N_RWLB<2>_XI814/MM9_g N_RBL<14>_XI814/MM9_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI814/MM6 N_XI814/NET08_XI814/MM6_d N_XI814/QB_XI814/MM6_g N_VDD_XI814/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI814/MM5 N_XI814/Q_XI814/MM5_d N_XI814/QB_XI814/MM5_g N_VDD_XI814/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI814/MM4 N_XI814/QB_XI814/MM4_d N_XI814/Q_XI814/MM4_g N_VDD_XI814/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI843/MM8 N_XI843/NET08_XI843/MM8_d N_RWL<3>_XI843/MM8_g N_RBL<1>_XI843/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI843/MM7 N_XI843/NET08_XI843/MM7_d N_XI843/QB_XI843/MM7_g N_GND_XI843/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI843/MM10 N_WBL<1>_XI843/MM10_d N_WWLB<3>_XI843/MM10_g N_XI843/Q_XI843/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI843/MM11 N_WBLB<1>_XI843/MM11_d N_WWLB<3>_XI843/MM11_g
+ N_XI843/QB_XI843/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI843/MM1 N_XI843/Q_XI843/MM1_d N_XI843/QB_XI843/MM1_g N_GND_XI843/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI843/MM0 N_XI843/QB_XI843/MM0_d N_XI843/Q_XI843/MM0_g N_GND_XI843/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI843/MM9 N_XI843/NET08_XI843/MM9_d N_RWLB<3>_XI843/MM9_g N_RBL<1>_XI843/MM9_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI843/MM6 N_XI843/NET08_XI843/MM6_d N_XI843/QB_XI843/MM6_g N_VDD_XI843/MM6_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI843/MM5 N_XI843/Q_XI843/MM5_d N_XI843/QB_XI843/MM5_g N_VDD_XI843/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI843/MM4 N_XI843/QB_XI843/MM4_d N_XI843/Q_XI843/MM4_g N_VDD_XI843/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI842/MM8 N_XI842/NET08_XI842/MM8_d N_RWL<3>_XI842/MM8_g N_RBL<2>_XI842/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI842/MM7 N_XI842/NET08_XI842/MM7_d N_XI842/QB_XI842/MM7_g N_GND_XI842/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI842/MM10 N_WBL<2>_XI842/MM10_d N_WWLB<3>_XI842/MM10_g N_XI842/Q_XI842/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI842/MM11 N_WBLB<2>_XI842/MM11_d N_WWLB<3>_XI842/MM11_g
+ N_XI842/QB_XI842/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI842/MM1 N_XI842/Q_XI842/MM1_d N_XI842/QB_XI842/MM1_g N_GND_XI842/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI842/MM0 N_XI842/QB_XI842/MM0_d N_XI842/Q_XI842/MM0_g N_GND_XI842/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI842/MM9 N_XI842/NET08_XI842/MM9_d N_RWLB<3>_XI842/MM9_g N_RBL<2>_XI842/MM9_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI842/MM6 N_XI842/NET08_XI842/MM6_d N_XI842/QB_XI842/MM6_g N_VDD_XI842/MM6_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI842/MM5 N_XI842/Q_XI842/MM5_d N_XI842/QB_XI842/MM5_g N_VDD_XI842/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI842/MM4 N_XI842/QB_XI842/MM4_d N_XI842/Q_XI842/MM4_g N_VDD_XI842/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI841/MM8 N_XI841/NET08_XI841/MM8_d N_RWL<3>_XI841/MM8_g N_RBL<3>_XI841/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI841/MM7 N_XI841/NET08_XI841/MM7_d N_XI841/QB_XI841/MM7_g N_GND_XI841/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI841/MM10 N_WBL<3>_XI841/MM10_d N_WWLB<3>_XI841/MM10_g N_XI841/Q_XI841/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI841/MM11 N_WBLB<3>_XI841/MM11_d N_WWLB<3>_XI841/MM11_g
+ N_XI841/QB_XI841/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI841/MM1 N_XI841/Q_XI841/MM1_d N_XI841/QB_XI841/MM1_g N_GND_XI841/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI841/MM0 N_XI841/QB_XI841/MM0_d N_XI841/Q_XI841/MM0_g N_GND_XI841/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI841/MM9 N_XI841/NET08_XI841/MM9_d N_RWLB<3>_XI841/MM9_g N_RBL<3>_XI841/MM9_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI841/MM6 N_XI841/NET08_XI841/MM6_d N_XI841/QB_XI841/MM6_g N_VDD_XI841/MM6_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI841/MM5 N_XI841/Q_XI841/MM5_d N_XI841/QB_XI841/MM5_g N_VDD_XI841/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI841/MM4 N_XI841/QB_XI841/MM4_d N_XI841/Q_XI841/MM4_g N_VDD_XI841/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI840/MM8 N_XI840/NET08_XI840/MM8_d N_RWL<3>_XI840/MM8_g N_RBL<4>_XI840/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI840/MM7 N_XI840/NET08_XI840/MM7_d N_XI840/QB_XI840/MM7_g N_GND_XI840/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI840/MM10 N_WBL<4>_XI840/MM10_d N_WWLB<3>_XI840/MM10_g N_XI840/Q_XI840/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI840/MM11 N_WBLB<4>_XI840/MM11_d N_WWLB<3>_XI840/MM11_g
+ N_XI840/QB_XI840/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI840/MM1 N_XI840/Q_XI840/MM1_d N_XI840/QB_XI840/MM1_g N_GND_XI840/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI840/MM0 N_XI840/QB_XI840/MM0_d N_XI840/Q_XI840/MM0_g N_GND_XI840/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI840/MM9 N_XI840/NET08_XI840/MM9_d N_RWLB<3>_XI840/MM9_g N_RBL<4>_XI840/MM9_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI840/MM6 N_XI840/NET08_XI840/MM6_d N_XI840/QB_XI840/MM6_g N_VDD_XI840/MM6_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI840/MM5 N_XI840/Q_XI840/MM5_d N_XI840/QB_XI840/MM5_g N_VDD_XI840/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI840/MM4 N_XI840/QB_XI840/MM4_d N_XI840/Q_XI840/MM4_g N_VDD_XI840/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1024/MM8 N_XI1024/NET08_XI1024/MM8_d N_RWL<15>_XI1024/MM8_g
+ N_RBL<12>_XI1024/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1024/MM7 N_XI1024/NET08_XI1024/MM7_d N_XI1024/QB_XI1024/MM7_g
+ N_GND_XI1024/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1024/MM10 N_WBL<12>_XI1024/MM10_d N_WWLB<15>_XI1024/MM10_g
+ N_XI1024/Q_XI1024/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1024/MM11 N_WBLB<12>_XI1024/MM11_d N_WWLB<15>_XI1024/MM11_g
+ N_XI1024/QB_XI1024/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1024/MM1 N_XI1024/Q_XI1024/MM1_d N_XI1024/QB_XI1024/MM1_g N_GND_XI1024/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1024/MM0 N_XI1024/QB_XI1024/MM0_d N_XI1024/Q_XI1024/MM0_g N_GND_XI1024/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1024/MM9 N_XI1024/NET08_XI1024/MM9_d N_RWLB<15>_XI1024/MM9_g
+ N_RBL<12>_XI1024/MM9_s N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1024/MM6 N_XI1024/NET08_XI1024/MM6_d N_XI1024/QB_XI1024/MM6_g
+ N_VDD_XI1024/MM6_s N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1024/MM5 N_XI1024/Q_XI1024/MM5_d N_XI1024/QB_XI1024/MM5_g N_VDD_XI1024/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1024/MM4 N_XI1024/QB_XI1024/MM4_d N_XI1024/Q_XI1024/MM4_g N_VDD_XI1024/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1003/MM8 N_XI1003/NET08_XI1003/MM8_d N_RWL<13>_XI1003/MM8_g
+ N_RBL<1>_XI1003/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1003/MM7 N_XI1003/NET08_XI1003/MM7_d N_XI1003/QB_XI1003/MM7_g
+ N_GND_XI1003/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1003/MM10 N_WBL<1>_XI1003/MM10_d N_WWLB<13>_XI1003/MM10_g
+ N_XI1003/Q_XI1003/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1003/MM11 N_WBLB<1>_XI1003/MM11_d N_WWLB<13>_XI1003/MM11_g
+ N_XI1003/QB_XI1003/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1003/MM1 N_XI1003/Q_XI1003/MM1_d N_XI1003/QB_XI1003/MM1_g N_GND_XI1003/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1003/MM0 N_XI1003/QB_XI1003/MM0_d N_XI1003/Q_XI1003/MM0_g N_GND_XI1003/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1003/MM9 N_XI1003/NET08_XI1003/MM9_d N_RWLB<13>_XI1003/MM9_g
+ N_RBL<1>_XI1003/MM9_s N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1003/MM6 N_XI1003/NET08_XI1003/MM6_d N_XI1003/QB_XI1003/MM6_g
+ N_VDD_XI1003/MM6_s N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1003/MM5 N_XI1003/Q_XI1003/MM5_d N_XI1003/QB_XI1003/MM5_g N_VDD_XI1003/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1003/MM4 N_XI1003/QB_XI1003/MM4_d N_XI1003/Q_XI1003/MM4_g N_VDD_XI1003/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI797/MM8 N_XI797/NET08_XI797/MM8_d N_RWL<0>_XI797/MM8_g N_RBL<0>_XI797/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI797/MM7 N_XI797/NET08_XI797/MM7_d N_XI797/QB_XI797/MM7_g N_GND_XI797/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI797/MM10 N_WBL<0>_XI797/MM10_d N_WWLB<0>_XI797/MM10_g N_XI797/Q_XI797/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI797/MM11 N_WBLB<0>_XI797/MM11_d N_WWLB<0>_XI797/MM11_g
+ N_XI797/QB_XI797/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI797/MM1 N_XI797/Q_XI797/MM1_d N_XI797/QB_XI797/MM1_g N_GND_XI797/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI797/MM0 N_XI797/QB_XI797/MM0_d N_XI797/Q_XI797/MM0_g N_GND_XI797/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI797/MM9 N_XI797/NET08_XI797/MM9_d N_RWLB<0>_XI797/MM9_g N_RBL<0>_XI797/MM9_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI797/MM6 N_XI797/NET08_XI797/MM6_d N_XI797/QB_XI797/MM6_g N_VDD_XI797/MM6_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI797/MM5 N_XI797/Q_XI797/MM5_d N_XI797/QB_XI797/MM5_g N_VDD_XI797/MM5_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI797/MM4 N_XI797/QB_XI797/MM4_d N_XI797/Q_XI797/MM4_g N_VDD_XI797/MM4_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI796/MM8 N_XI796/NET08_XI796/MM8_d N_RWL<0>_XI796/MM8_g N_RBL<1>_XI796/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI796/MM7 N_XI796/NET08_XI796/MM7_d N_XI796/QB_XI796/MM7_g N_GND_XI796/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI796/MM10 N_WBL<1>_XI796/MM10_d N_WWLB<0>_XI796/MM10_g N_XI796/Q_XI796/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI796/MM11 N_WBLB<1>_XI796/MM11_d N_WWLB<0>_XI796/MM11_g
+ N_XI796/QB_XI796/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI796/MM1 N_XI796/Q_XI796/MM1_d N_XI796/QB_XI796/MM1_g N_GND_XI796/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI796/MM0 N_XI796/QB_XI796/MM0_d N_XI796/Q_XI796/MM0_g N_GND_XI796/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI796/MM9 N_XI796/NET08_XI796/MM9_d N_RWLB<0>_XI796/MM9_g N_RBL<1>_XI796/MM9_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI796/MM6 N_XI796/NET08_XI796/MM6_d N_XI796/QB_XI796/MM6_g N_VDD_XI796/MM6_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI796/MM5 N_XI796/Q_XI796/MM5_d N_XI796/QB_XI796/MM5_g N_VDD_XI796/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI796/MM4 N_XI796/QB_XI796/MM4_d N_XI796/Q_XI796/MM4_g N_VDD_XI796/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI795/MM8 N_XI795/NET08_XI795/MM8_d N_RWL<0>_XI795/MM8_g N_RBL<2>_XI795/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI795/MM7 N_XI795/NET08_XI795/MM7_d N_XI795/QB_XI795/MM7_g N_GND_XI795/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI795/MM10 N_WBL<2>_XI795/MM10_d N_WWLB<0>_XI795/MM10_g N_XI795/Q_XI795/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI795/MM11 N_WBLB<2>_XI795/MM11_d N_WWLB<0>_XI795/MM11_g
+ N_XI795/QB_XI795/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI795/MM1 N_XI795/Q_XI795/MM1_d N_XI795/QB_XI795/MM1_g N_GND_XI795/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI795/MM0 N_XI795/QB_XI795/MM0_d N_XI795/Q_XI795/MM0_g N_GND_XI795/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI795/MM9 N_XI795/NET08_XI795/MM9_d N_RWLB<0>_XI795/MM9_g N_RBL<2>_XI795/MM9_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI795/MM6 N_XI795/NET08_XI795/MM6_d N_XI795/QB_XI795/MM6_g N_VDD_XI795/MM6_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI795/MM5 N_XI795/Q_XI795/MM5_d N_XI795/QB_XI795/MM5_g N_VDD_XI795/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI795/MM4 N_XI795/QB_XI795/MM4_d N_XI795/Q_XI795/MM4_g N_VDD_XI795/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI788/MM8 N_XI788/NET08_XI788/MM8_d N_RWL<0>_XI788/MM8_g N_RBL<9>_XI788/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI788/MM7 N_XI788/NET08_XI788/MM7_d N_XI788/QB_XI788/MM7_g N_GND_XI788/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI788/MM10 N_WBL<9>_XI788/MM10_d N_WWLB<0>_XI788/MM10_g N_XI788/Q_XI788/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI788/MM11 N_WBLB<9>_XI788/MM11_d N_WWLB<0>_XI788/MM11_g
+ N_XI788/QB_XI788/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI788/MM1 N_XI788/Q_XI788/MM1_d N_XI788/QB_XI788/MM1_g N_GND_XI788/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI788/MM0 N_XI788/QB_XI788/MM0_d N_XI788/Q_XI788/MM0_g N_GND_XI788/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI788/MM9 N_XI788/NET08_XI788/MM9_d N_RWLB<0>_XI788/MM9_g N_RBL<9>_XI788/MM9_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI788/MM6 N_XI788/NET08_XI788/MM6_d N_XI788/QB_XI788/MM6_g N_VDD_XI788/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI788/MM5 N_XI788/Q_XI788/MM5_d N_XI788/QB_XI788/MM5_g N_VDD_XI788/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI788/MM4 N_XI788/QB_XI788/MM4_d N_XI788/Q_XI788/MM4_g N_VDD_XI788/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI787/MM8 N_XI787/NET08_XI787/MM8_d N_RWL<0>_XI787/MM8_g N_RBL<10>_XI787/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI787/MM7 N_XI787/NET08_XI787/MM7_d N_XI787/QB_XI787/MM7_g N_GND_XI787/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI787/MM10 N_WBL<10>_XI787/MM10_d N_WWLB<0>_XI787/MM10_g N_XI787/Q_XI787/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI787/MM11 N_WBLB<10>_XI787/MM11_d N_WWLB<0>_XI787/MM11_g
+ N_XI787/QB_XI787/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI787/MM1 N_XI787/Q_XI787/MM1_d N_XI787/QB_XI787/MM1_g N_GND_XI787/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI787/MM0 N_XI787/QB_XI787/MM0_d N_XI787/Q_XI787/MM0_g N_GND_XI787/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI787/MM9 N_XI787/NET08_XI787/MM9_d N_RWLB<0>_XI787/MM9_g N_RBL<10>_XI787/MM9_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI787/MM6 N_XI787/NET08_XI787/MM6_d N_XI787/QB_XI787/MM6_g N_VDD_XI787/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI787/MM5 N_XI787/Q_XI787/MM5_d N_XI787/QB_XI787/MM5_g N_VDD_XI787/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI787/MM4 N_XI787/QB_XI787/MM4_d N_XI787/Q_XI787/MM4_g N_VDD_XI787/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI786/MM8 N_XI786/NET08_XI786/MM8_d N_RWL<0>_XI786/MM8_g N_RBL<11>_XI786/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI786/MM7 N_XI786/NET08_XI786/MM7_d N_XI786/QB_XI786/MM7_g N_GND_XI786/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI786/MM10 N_WBL<11>_XI786/MM10_d N_WWLB<0>_XI786/MM10_g N_XI786/Q_XI786/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI786/MM11 N_WBLB<11>_XI786/MM11_d N_WWLB<0>_XI786/MM11_g
+ N_XI786/QB_XI786/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI786/MM1 N_XI786/Q_XI786/MM1_d N_XI786/QB_XI786/MM1_g N_GND_XI786/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI786/MM0 N_XI786/QB_XI786/MM0_d N_XI786/Q_XI786/MM0_g N_GND_XI786/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI786/MM9 N_XI786/NET08_XI786/MM9_d N_RWLB<0>_XI786/MM9_g N_RBL<11>_XI786/MM9_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI786/MM6 N_XI786/NET08_XI786/MM6_d N_XI786/QB_XI786/MM6_g N_VDD_XI786/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI786/MM5 N_XI786/Q_XI786/MM5_d N_XI786/QB_XI786/MM5_g N_VDD_XI786/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI786/MM4 N_XI786/QB_XI786/MM4_d N_XI786/Q_XI786/MM4_g N_VDD_XI786/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI813/MM8 N_XI813/NET08_XI813/MM8_d N_RWL<1>_XI813/MM8_g N_RBL<15>_XI813/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI813/MM7 N_XI813/NET08_XI813/MM7_d N_XI813/QB_XI813/MM7_g N_GND_XI813/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI813/MM10 N_WBL<15>_XI813/MM10_d N_WWLB<1>_XI813/MM10_g N_XI813/Q_XI813/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI813/MM11 N_WBLB<15>_XI813/MM11_d N_WWLB<1>_XI813/MM11_g
+ N_XI813/QB_XI813/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI813/MM1 N_XI813/Q_XI813/MM1_d N_XI813/QB_XI813/MM1_g N_GND_XI813/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI813/MM0 N_XI813/QB_XI813/MM0_d N_XI813/Q_XI813/MM0_g N_GND_XI813/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI813/MM9 N_XI813/NET08_XI813/MM9_d N_RWLB<1>_XI813/MM9_g N_RBL<15>_XI813/MM9_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI813/MM6 N_XI813/NET08_XI813/MM6_d N_XI813/QB_XI813/MM6_g N_VDD_XI813/MM6_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI813/MM5 N_XI813/Q_XI813/MM5_d N_XI813/QB_XI813/MM5_g N_VDD_XI813/MM5_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI813/MM4 N_XI813/QB_XI813/MM4_d N_XI813/Q_XI813/MM4_g N_VDD_XI813/MM4_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI812/MM8 N_XI812/NET08_XI812/MM8_d N_RWL<1>_XI812/MM8_g N_RBL<0>_XI812/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI812/MM7 N_XI812/NET08_XI812/MM7_d N_XI812/QB_XI812/MM7_g N_GND_XI812/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI812/MM10 N_WBL<0>_XI812/MM10_d N_WWLB<1>_XI812/MM10_g N_XI812/Q_XI812/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI812/MM11 N_WBLB<0>_XI812/MM11_d N_WWLB<1>_XI812/MM11_g
+ N_XI812/QB_XI812/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI812/MM1 N_XI812/Q_XI812/MM1_d N_XI812/QB_XI812/MM1_g N_GND_XI812/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI812/MM0 N_XI812/QB_XI812/MM0_d N_XI812/Q_XI812/MM0_g N_GND_XI812/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI812/MM9 N_XI812/NET08_XI812/MM9_d N_RWLB<1>_XI812/MM9_g N_RBL<0>_XI812/MM9_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI812/MM6 N_XI812/NET08_XI812/MM6_d N_XI812/QB_XI812/MM6_g N_VDD_XI812/MM6_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI812/MM5 N_XI812/Q_XI812/MM5_d N_XI812/QB_XI812/MM5_g N_VDD_XI812/MM5_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI812/MM4 N_XI812/QB_XI812/MM4_d N_XI812/Q_XI812/MM4_g N_VDD_XI812/MM4_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI811/MM8 N_XI811/NET08_XI811/MM8_d N_RWL<1>_XI811/MM8_g N_RBL<1>_XI811/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI811/MM7 N_XI811/NET08_XI811/MM7_d N_XI811/QB_XI811/MM7_g N_GND_XI811/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI811/MM10 N_WBL<1>_XI811/MM10_d N_WWLB<1>_XI811/MM10_g N_XI811/Q_XI811/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI811/MM11 N_WBLB<1>_XI811/MM11_d N_WWLB<1>_XI811/MM11_g
+ N_XI811/QB_XI811/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI811/MM1 N_XI811/Q_XI811/MM1_d N_XI811/QB_XI811/MM1_g N_GND_XI811/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI811/MM0 N_XI811/QB_XI811/MM0_d N_XI811/Q_XI811/MM0_g N_GND_XI811/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI811/MM9 N_XI811/NET08_XI811/MM9_d N_RWLB<1>_XI811/MM9_g N_RBL<1>_XI811/MM9_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI811/MM6 N_XI811/NET08_XI811/MM6_d N_XI811/QB_XI811/MM6_g N_VDD_XI811/MM6_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI811/MM5 N_XI811/Q_XI811/MM5_d N_XI811/QB_XI811/MM5_g N_VDD_XI811/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI811/MM4 N_XI811/QB_XI811/MM4_d N_XI811/Q_XI811/MM4_g N_VDD_XI811/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI810/MM8 N_XI810/NET08_XI810/MM8_d N_RWL<1>_XI810/MM8_g N_RBL<2>_XI810/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI810/MM7 N_XI810/NET08_XI810/MM7_d N_XI810/QB_XI810/MM7_g N_GND_XI810/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI810/MM10 N_WBL<2>_XI810/MM10_d N_WWLB<1>_XI810/MM10_g N_XI810/Q_XI810/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI810/MM11 N_WBLB<2>_XI810/MM11_d N_WWLB<1>_XI810/MM11_g
+ N_XI810/QB_XI810/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI810/MM1 N_XI810/Q_XI810/MM1_d N_XI810/QB_XI810/MM1_g N_GND_XI810/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI810/MM0 N_XI810/QB_XI810/MM0_d N_XI810/Q_XI810/MM0_g N_GND_XI810/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI810/MM9 N_XI810/NET08_XI810/MM9_d N_RWLB<1>_XI810/MM9_g N_RBL<2>_XI810/MM9_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI810/MM6 N_XI810/NET08_XI810/MM6_d N_XI810/QB_XI810/MM6_g N_VDD_XI810/MM6_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI810/MM5 N_XI810/Q_XI810/MM5_d N_XI810/QB_XI810/MM5_g N_VDD_XI810/MM5_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI810/MM4 N_XI810/QB_XI810/MM4_d N_XI810/Q_XI810/MM4_g N_VDD_XI810/MM4_s
+ N_VDD_XI1034/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI809/MM8 N_XI809/NET08_XI809/MM8_d N_RWL<1>_XI809/MM8_g N_RBL<3>_XI809/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI809/MM7 N_XI809/NET08_XI809/MM7_d N_XI809/QB_XI809/MM7_g N_GND_XI809/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI809/MM10 N_WBL<3>_XI809/MM10_d N_WWLB<1>_XI809/MM10_g N_XI809/Q_XI809/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI809/MM11 N_WBLB<3>_XI809/MM11_d N_WWLB<1>_XI809/MM11_g
+ N_XI809/QB_XI809/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI809/MM1 N_XI809/Q_XI809/MM1_d N_XI809/QB_XI809/MM1_g N_GND_XI809/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI809/MM0 N_XI809/QB_XI809/MM0_d N_XI809/Q_XI809/MM0_g N_GND_XI809/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI809/MM9 N_XI809/NET08_XI809/MM9_d N_RWLB<1>_XI809/MM9_g N_RBL<3>_XI809/MM9_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI809/MM6 N_XI809/NET08_XI809/MM6_d N_XI809/QB_XI809/MM6_g N_VDD_XI809/MM6_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI809/MM5 N_XI809/Q_XI809/MM5_d N_XI809/QB_XI809/MM5_g N_VDD_XI809/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI809/MM4 N_XI809/QB_XI809/MM4_d N_XI809/Q_XI809/MM4_g N_VDD_XI809/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI808/MM8 N_XI808/NET08_XI808/MM8_d N_RWL<1>_XI808/MM8_g N_RBL<4>_XI808/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI808/MM7 N_XI808/NET08_XI808/MM7_d N_XI808/QB_XI808/MM7_g N_GND_XI808/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI808/MM10 N_WBL<4>_XI808/MM10_d N_WWLB<1>_XI808/MM10_g N_XI808/Q_XI808/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI808/MM11 N_WBLB<4>_XI808/MM11_d N_WWLB<1>_XI808/MM11_g
+ N_XI808/QB_XI808/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI808/MM1 N_XI808/Q_XI808/MM1_d N_XI808/QB_XI808/MM1_g N_GND_XI808/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI808/MM0 N_XI808/QB_XI808/MM0_d N_XI808/Q_XI808/MM0_g N_GND_XI808/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI808/MM9 N_XI808/NET08_XI808/MM9_d N_RWLB<1>_XI808/MM9_g N_RBL<4>_XI808/MM9_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI808/MM6 N_XI808/NET08_XI808/MM6_d N_XI808/QB_XI808/MM6_g N_VDD_XI808/MM6_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI808/MM5 N_XI808/Q_XI808/MM5_d N_XI808/QB_XI808/MM5_g N_VDD_XI808/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI808/MM4 N_XI808/QB_XI808/MM4_d N_XI808/Q_XI808/MM4_g N_VDD_XI808/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI839/MM8 N_XI839/NET08_XI839/MM8_d N_RWL<3>_XI839/MM8_g N_RBL<5>_XI839/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI839/MM7 N_XI839/NET08_XI839/MM7_d N_XI839/QB_XI839/MM7_g N_GND_XI839/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI839/MM10 N_WBL<5>_XI839/MM10_d N_WWLB<3>_XI839/MM10_g N_XI839/Q_XI839/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI839/MM11 N_WBLB<5>_XI839/MM11_d N_WWLB<3>_XI839/MM11_g
+ N_XI839/QB_XI839/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI839/MM1 N_XI839/Q_XI839/MM1_d N_XI839/QB_XI839/MM1_g N_GND_XI839/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI839/MM0 N_XI839/QB_XI839/MM0_d N_XI839/Q_XI839/MM0_g N_GND_XI839/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI839/MM9 N_XI839/NET08_XI839/MM9_d N_RWLB<3>_XI839/MM9_g N_RBL<5>_XI839/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI839/MM6 N_XI839/NET08_XI839/MM6_d N_XI839/QB_XI839/MM6_g N_VDD_XI839/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI839/MM5 N_XI839/Q_XI839/MM5_d N_XI839/QB_XI839/MM5_g N_VDD_XI839/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI839/MM4 N_XI839/QB_XI839/MM4_d N_XI839/Q_XI839/MM4_g N_VDD_XI839/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI838/MM8 N_XI838/NET08_XI838/MM8_d N_RWL<3>_XI838/MM8_g N_RBL<6>_XI838/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI838/MM7 N_XI838/NET08_XI838/MM7_d N_XI838/QB_XI838/MM7_g N_GND_XI838/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI838/MM10 N_WBL<6>_XI838/MM10_d N_WWLB<3>_XI838/MM10_g N_XI838/Q_XI838/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI838/MM11 N_WBLB<6>_XI838/MM11_d N_WWLB<3>_XI838/MM11_g
+ N_XI838/QB_XI838/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI838/MM1 N_XI838/Q_XI838/MM1_d N_XI838/QB_XI838/MM1_g N_GND_XI838/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI838/MM0 N_XI838/QB_XI838/MM0_d N_XI838/Q_XI838/MM0_g N_GND_XI838/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI838/MM9 N_XI838/NET08_XI838/MM9_d N_RWLB<3>_XI838/MM9_g N_RBL<6>_XI838/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI838/MM6 N_XI838/NET08_XI838/MM6_d N_XI838/QB_XI838/MM6_g N_VDD_XI838/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI838/MM5 N_XI838/Q_XI838/MM5_d N_XI838/QB_XI838/MM5_g N_VDD_XI838/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI838/MM4 N_XI838/QB_XI838/MM4_d N_XI838/Q_XI838/MM4_g N_VDD_XI838/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI837/MM8 N_XI837/NET08_XI837/MM8_d N_RWL<3>_XI837/MM8_g N_RBL<7>_XI837/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI837/MM7 N_XI837/NET08_XI837/MM7_d N_XI837/QB_XI837/MM7_g N_GND_XI837/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI837/MM10 N_WBL<7>_XI837/MM10_d N_WWLB<3>_XI837/MM10_g N_XI837/Q_XI837/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI837/MM11 N_WBLB<7>_XI837/MM11_d N_WWLB<3>_XI837/MM11_g
+ N_XI837/QB_XI837/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI837/MM1 N_XI837/Q_XI837/MM1_d N_XI837/QB_XI837/MM1_g N_GND_XI837/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI837/MM0 N_XI837/QB_XI837/MM0_d N_XI837/Q_XI837/MM0_g N_GND_XI837/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI837/MM9 N_XI837/NET08_XI837/MM9_d N_RWLB<3>_XI837/MM9_g N_RBL<7>_XI837/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI837/MM6 N_XI837/NET08_XI837/MM6_d N_XI837/QB_XI837/MM6_g N_VDD_XI837/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI837/MM5 N_XI837/Q_XI837/MM5_d N_XI837/QB_XI837/MM5_g N_VDD_XI837/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI837/MM4 N_XI837/QB_XI837/MM4_d N_XI837/Q_XI837/MM4_g N_VDD_XI837/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI836/MM8 N_XI836/NET08_XI836/MM8_d N_RWL<3>_XI836/MM8_g N_RBL<8>_XI836/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI836/MM7 N_XI836/NET08_XI836/MM7_d N_XI836/QB_XI836/MM7_g N_GND_XI836/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI836/MM10 N_WBL<8>_XI836/MM10_d N_WWLB<3>_XI836/MM10_g N_XI836/Q_XI836/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI836/MM11 N_WBLB<8>_XI836/MM11_d N_WWLB<3>_XI836/MM11_g
+ N_XI836/QB_XI836/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI836/MM1 N_XI836/Q_XI836/MM1_d N_XI836/QB_XI836/MM1_g N_GND_XI836/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI836/MM0 N_XI836/QB_XI836/MM0_d N_XI836/Q_XI836/MM0_g N_GND_XI836/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI836/MM9 N_XI836/NET08_XI836/MM9_d N_RWLB<3>_XI836/MM9_g N_RBL<8>_XI836/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI836/MM6 N_XI836/NET08_XI836/MM6_d N_XI836/QB_XI836/MM6_g N_VDD_XI836/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI836/MM5 N_XI836/Q_XI836/MM5_d N_XI836/QB_XI836/MM5_g N_VDD_XI836/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI836/MM4 N_XI836/QB_XI836/MM4_d N_XI836/Q_XI836/MM4_g N_VDD_XI836/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1023/MM8 N_XI1023/NET08_XI1023/MM8_d N_RWL<15>_XI1023/MM8_g
+ N_RBL<13>_XI1023/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1023/MM7 N_XI1023/NET08_XI1023/MM7_d N_XI1023/QB_XI1023/MM7_g
+ N_GND_XI1023/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1023/MM10 N_WBL<13>_XI1023/MM10_d N_WWLB<15>_XI1023/MM10_g
+ N_XI1023/Q_XI1023/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1023/MM11 N_WBLB<13>_XI1023/MM11_d N_WWLB<15>_XI1023/MM11_g
+ N_XI1023/QB_XI1023/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1023/MM1 N_XI1023/Q_XI1023/MM1_d N_XI1023/QB_XI1023/MM1_g N_GND_XI1023/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1023/MM0 N_XI1023/QB_XI1023/MM0_d N_XI1023/Q_XI1023/MM0_g N_GND_XI1023/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1023/MM9 N_XI1023/NET08_XI1023/MM9_d N_RWLB<15>_XI1023/MM9_g
+ N_RBL<13>_XI1023/MM9_s N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1023/MM6 N_XI1023/NET08_XI1023/MM6_d N_XI1023/QB_XI1023/MM6_g
+ N_VDD_XI1023/MM6_s N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1023/MM5 N_XI1023/Q_XI1023/MM5_d N_XI1023/QB_XI1023/MM5_g N_VDD_XI1023/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1023/MM4 N_XI1023/QB_XI1023/MM4_d N_XI1023/Q_XI1023/MM4_g N_VDD_XI1023/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1004/MM8 N_XI1004/NET08_XI1004/MM8_d N_RWL<13>_XI1004/MM8_g
+ N_RBL<0>_XI1004/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1004/MM7 N_XI1004/NET08_XI1004/MM7_d N_XI1004/QB_XI1004/MM7_g
+ N_GND_XI1004/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1004/MM10 N_WBL<0>_XI1004/MM10_d N_WWLB<13>_XI1004/MM10_g
+ N_XI1004/Q_XI1004/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1004/MM11 N_WBLB<0>_XI1004/MM11_d N_WWLB<13>_XI1004/MM11_g
+ N_XI1004/QB_XI1004/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1004/MM1 N_XI1004/Q_XI1004/MM1_d N_XI1004/QB_XI1004/MM1_g N_GND_XI1004/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1004/MM0 N_XI1004/QB_XI1004/MM0_d N_XI1004/Q_XI1004/MM0_g N_GND_XI1004/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1004/MM9 N_XI1004/NET08_XI1004/MM9_d N_RWLB<13>_XI1004/MM9_g
+ N_RBL<0>_XI1004/MM9_s N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1004/MM6 N_XI1004/NET08_XI1004/MM6_d N_XI1004/QB_XI1004/MM6_g
+ N_VDD_XI1004/MM6_s N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1004/MM5 N_XI1004/Q_XI1004/MM5_d N_XI1004/QB_XI1004/MM5_g N_VDD_XI1004/MM5_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1004/MM4 N_XI1004/QB_XI1004/MM4_d N_XI1004/Q_XI1004/MM4_g N_VDD_XI1004/MM4_s
+ N_VDD_XI1036/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI793/MM8 N_XI793/NET08_XI793/MM8_d N_RWL<0>_XI793/MM8_g N_RBL<4>_XI793/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI793/MM7 N_XI793/NET08_XI793/MM7_d N_XI793/QB_XI793/MM7_g N_GND_XI793/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI793/MM10 N_WBL<4>_XI793/MM10_d N_WWLB<0>_XI793/MM10_g N_XI793/Q_XI793/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI793/MM11 N_WBLB<4>_XI793/MM11_d N_WWLB<0>_XI793/MM11_g
+ N_XI793/QB_XI793/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI793/MM1 N_XI793/Q_XI793/MM1_d N_XI793/QB_XI793/MM1_g N_GND_XI793/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI793/MM0 N_XI793/QB_XI793/MM0_d N_XI793/Q_XI793/MM0_g N_GND_XI793/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI793/MM9 N_XI793/NET08_XI793/MM9_d N_RWLB<0>_XI793/MM9_g N_RBL<4>_XI793/MM9_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI793/MM6 N_XI793/NET08_XI793/MM6_d N_XI793/QB_XI793/MM6_g N_VDD_XI793/MM6_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI793/MM5 N_XI793/Q_XI793/MM5_d N_XI793/QB_XI793/MM5_g N_VDD_XI793/MM5_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI793/MM4 N_XI793/QB_XI793/MM4_d N_XI793/Q_XI793/MM4_g N_VDD_XI793/MM4_s
+ N_VDD_XI1032/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI792/MM8 N_XI792/NET08_XI792/MM8_d N_RWL<0>_XI792/MM8_g N_RBL<5>_XI792/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI792/MM7 N_XI792/NET08_XI792/MM7_d N_XI792/QB_XI792/MM7_g N_GND_XI792/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI792/MM10 N_WBL<5>_XI792/MM10_d N_WWLB<0>_XI792/MM10_g N_XI792/Q_XI792/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI792/MM11 N_WBLB<5>_XI792/MM11_d N_WWLB<0>_XI792/MM11_g
+ N_XI792/QB_XI792/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI792/MM1 N_XI792/Q_XI792/MM1_d N_XI792/QB_XI792/MM1_g N_GND_XI792/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI792/MM0 N_XI792/QB_XI792/MM0_d N_XI792/Q_XI792/MM0_g N_GND_XI792/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI792/MM9 N_XI792/NET08_XI792/MM9_d N_RWLB<0>_XI792/MM9_g N_RBL<5>_XI792/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI792/MM6 N_XI792/NET08_XI792/MM6_d N_XI792/QB_XI792/MM6_g N_VDD_XI792/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI792/MM5 N_XI792/Q_XI792/MM5_d N_XI792/QB_XI792/MM5_g N_VDD_XI792/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI792/MM4 N_XI792/QB_XI792/MM4_d N_XI792/Q_XI792/MM4_g N_VDD_XI792/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI784/MM8 N_XI784/NET08_XI784/MM8_d N_RWL<0>_XI784/MM8_g N_RBL<13>_XI784/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI784/MM7 N_XI784/NET08_XI784/MM7_d N_XI784/QB_XI784/MM7_g N_GND_XI784/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI784/MM10 N_WBL<13>_XI784/MM10_d N_WWLB<0>_XI784/MM10_g N_XI784/Q_XI784/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI784/MM11 N_WBLB<13>_XI784/MM11_d N_WWLB<0>_XI784/MM11_g
+ N_XI784/QB_XI784/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI784/MM1 N_XI784/Q_XI784/MM1_d N_XI784/QB_XI784/MM1_g N_GND_XI784/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI784/MM0 N_XI784/QB_XI784/MM0_d N_XI784/Q_XI784/MM0_g N_GND_XI784/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI784/MM9 N_XI784/NET08_XI784/MM9_d N_RWLB<0>_XI784/MM9_g N_RBL<13>_XI784/MM9_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI784/MM6 N_XI784/NET08_XI784/MM6_d N_XI784/QB_XI784/MM6_g N_VDD_XI784/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI784/MM5 N_XI784/Q_XI784/MM5_d N_XI784/QB_XI784/MM5_g N_VDD_XI784/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI784/MM4 N_XI784/QB_XI784/MM4_d N_XI784/Q_XI784/MM4_g N_VDD_XI784/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI783/MM8 N_XI783/NET08_XI783/MM8_d N_RWL<0>_XI783/MM8_g N_RBL<14>_XI783/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI783/MM7 N_XI783/NET08_XI783/MM7_d N_XI783/QB_XI783/MM7_g N_GND_XI783/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI783/MM10 N_WBL<14>_XI783/MM10_d N_WWLB<0>_XI783/MM10_g N_XI783/Q_XI783/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI783/MM11 N_WBLB<14>_XI783/MM11_d N_WWLB<0>_XI783/MM11_g
+ N_XI783/QB_XI783/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI783/MM1 N_XI783/Q_XI783/MM1_d N_XI783/QB_XI783/MM1_g N_GND_XI783/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI783/MM0 N_XI783/QB_XI783/MM0_d N_XI783/Q_XI783/MM0_g N_GND_XI783/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI783/MM9 N_XI783/NET08_XI783/MM9_d N_RWLB<0>_XI783/MM9_g N_RBL<14>_XI783/MM9_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI783/MM6 N_XI783/NET08_XI783/MM6_d N_XI783/QB_XI783/MM6_g N_VDD_XI783/MM6_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI783/MM5 N_XI783/Q_XI783/MM5_d N_XI783/QB_XI783/MM5_g N_VDD_XI783/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI783/MM4 N_XI783/QB_XI783/MM4_d N_XI783/Q_XI783/MM4_g N_VDD_XI783/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI782/MM8 N_XI782/NET08_XI782/MM8_d N_RWL<0>_XI782/MM8_g N_RBL<15>_XI782/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI782/MM7 N_XI782/NET08_XI782/MM7_d N_XI782/QB_XI782/MM7_g N_GND_XI782/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI782/MM10 N_WBL<15>_XI782/MM10_d N_WWLB<0>_XI782/MM10_g N_XI782/Q_XI782/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI782/MM11 N_WBLB<15>_XI782/MM11_d N_WWLB<0>_XI782/MM11_g
+ N_XI782/QB_XI782/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI782/MM1 N_XI782/Q_XI782/MM1_d N_XI782/QB_XI782/MM1_g N_GND_XI782/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI782/MM0 N_XI782/QB_XI782/MM0_d N_XI782/Q_XI782/MM0_g N_GND_XI782/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI782/MM9 N_XI782/NET08_XI782/MM9_d N_RWLB<0>_XI782/MM9_g N_RBL<15>_XI782/MM9_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI782/MM6 N_XI782/NET08_XI782/MM6_d N_XI782/QB_XI782/MM6_g N_VDD_XI782/MM6_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI782/MM5 N_XI782/Q_XI782/MM5_d N_XI782/QB_XI782/MM5_g N_VDD_XI782/MM5_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI782/MM4 N_XI782/QB_XI782/MM4_d N_XI782/Q_XI782/MM4_g N_VDD_XI782/MM4_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI785/MM8 N_XI785/NET08_XI785/MM8_d N_RWL<0>_XI785/MM8_g N_RBL<12>_XI785/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI785/MM7 N_XI785/NET08_XI785/MM7_d N_XI785/QB_XI785/MM7_g N_GND_XI785/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI785/MM10 N_WBL<12>_XI785/MM10_d N_WWLB<0>_XI785/MM10_g N_XI785/Q_XI785/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI785/MM11 N_WBLB<12>_XI785/MM11_d N_WWLB<0>_XI785/MM11_g
+ N_XI785/QB_XI785/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI785/MM1 N_XI785/Q_XI785/MM1_d N_XI785/QB_XI785/MM1_g N_GND_XI785/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI785/MM0 N_XI785/QB_XI785/MM0_d N_XI785/Q_XI785/MM0_g N_GND_XI785/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI785/MM9 N_XI785/NET08_XI785/MM9_d N_RWLB<0>_XI785/MM9_g N_RBL<12>_XI785/MM9_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI785/MM6 N_XI785/NET08_XI785/MM6_d N_XI785/QB_XI785/MM6_g N_VDD_XI785/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI785/MM5 N_XI785/Q_XI785/MM5_d N_XI785/QB_XI785/MM5_g N_VDD_XI785/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI785/MM4 N_XI785/QB_XI785/MM4_d N_XI785/Q_XI785/MM4_g N_VDD_XI785/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI806/MM8 N_XI806/NET08_XI806/MM8_d N_RWL<1>_XI806/MM8_g N_RBL<6>_XI806/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI806/MM7 N_XI806/NET08_XI806/MM7_d N_XI806/QB_XI806/MM7_g N_GND_XI806/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI806/MM10 N_WBL<6>_XI806/MM10_d N_WWLB<1>_XI806/MM10_g N_XI806/Q_XI806/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI806/MM11 N_WBLB<6>_XI806/MM11_d N_WWLB<1>_XI806/MM11_g
+ N_XI806/QB_XI806/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI806/MM1 N_XI806/Q_XI806/MM1_d N_XI806/QB_XI806/MM1_g N_GND_XI806/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI806/MM0 N_XI806/QB_XI806/MM0_d N_XI806/Q_XI806/MM0_g N_GND_XI806/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI806/MM9 N_XI806/NET08_XI806/MM9_d N_RWLB<1>_XI806/MM9_g N_RBL<6>_XI806/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI806/MM6 N_XI806/NET08_XI806/MM6_d N_XI806/QB_XI806/MM6_g N_VDD_XI806/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI806/MM5 N_XI806/Q_XI806/MM5_d N_XI806/QB_XI806/MM5_g N_VDD_XI806/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI806/MM4 N_XI806/QB_XI806/MM4_d N_XI806/Q_XI806/MM4_g N_VDD_XI806/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI805/MM8 N_XI805/NET08_XI805/MM8_d N_RWL<1>_XI805/MM8_g N_RBL<7>_XI805/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI805/MM7 N_XI805/NET08_XI805/MM7_d N_XI805/QB_XI805/MM7_g N_GND_XI805/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI805/MM10 N_WBL<7>_XI805/MM10_d N_WWLB<1>_XI805/MM10_g N_XI805/Q_XI805/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI805/MM11 N_WBLB<7>_XI805/MM11_d N_WWLB<1>_XI805/MM11_g
+ N_XI805/QB_XI805/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI805/MM1 N_XI805/Q_XI805/MM1_d N_XI805/QB_XI805/MM1_g N_GND_XI805/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI805/MM0 N_XI805/QB_XI805/MM0_d N_XI805/Q_XI805/MM0_g N_GND_XI805/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI805/MM9 N_XI805/NET08_XI805/MM9_d N_RWLB<1>_XI805/MM9_g N_RBL<7>_XI805/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI805/MM6 N_XI805/NET08_XI805/MM6_d N_XI805/QB_XI805/MM6_g N_VDD_XI805/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI805/MM5 N_XI805/Q_XI805/MM5_d N_XI805/QB_XI805/MM5_g N_VDD_XI805/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI805/MM4 N_XI805/QB_XI805/MM4_d N_XI805/Q_XI805/MM4_g N_VDD_XI805/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI804/MM8 N_XI804/NET08_XI804/MM8_d N_RWL<1>_XI804/MM8_g N_RBL<8>_XI804/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI804/MM7 N_XI804/NET08_XI804/MM7_d N_XI804/QB_XI804/MM7_g N_GND_XI804/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI804/MM10 N_WBL<8>_XI804/MM10_d N_WWLB<1>_XI804/MM10_g N_XI804/Q_XI804/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI804/MM11 N_WBLB<8>_XI804/MM11_d N_WWLB<1>_XI804/MM11_g
+ N_XI804/QB_XI804/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI804/MM1 N_XI804/Q_XI804/MM1_d N_XI804/QB_XI804/MM1_g N_GND_XI804/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI804/MM0 N_XI804/QB_XI804/MM0_d N_XI804/Q_XI804/MM0_g N_GND_XI804/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI804/MM9 N_XI804/NET08_XI804/MM9_d N_RWLB<1>_XI804/MM9_g N_RBL<8>_XI804/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI804/MM6 N_XI804/NET08_XI804/MM6_d N_XI804/QB_XI804/MM6_g N_VDD_XI804/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI804/MM5 N_XI804/Q_XI804/MM5_d N_XI804/QB_XI804/MM5_g N_VDD_XI804/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI804/MM4 N_XI804/QB_XI804/MM4_d N_XI804/Q_XI804/MM4_g N_VDD_XI804/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI803/MM8 N_XI803/NET08_XI803/MM8_d N_RWL<1>_XI803/MM8_g N_RBL<9>_XI803/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI803/MM7 N_XI803/NET08_XI803/MM7_d N_XI803/QB_XI803/MM7_g N_GND_XI803/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI803/MM10 N_WBL<9>_XI803/MM10_d N_WWLB<1>_XI803/MM10_g N_XI803/Q_XI803/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI803/MM11 N_WBLB<9>_XI803/MM11_d N_WWLB<1>_XI803/MM11_g
+ N_XI803/QB_XI803/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI803/MM1 N_XI803/Q_XI803/MM1_d N_XI803/QB_XI803/MM1_g N_GND_XI803/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI803/MM0 N_XI803/QB_XI803/MM0_d N_XI803/Q_XI803/MM0_g N_GND_XI803/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI803/MM9 N_XI803/NET08_XI803/MM9_d N_RWLB<1>_XI803/MM9_g N_RBL<9>_XI803/MM9_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI803/MM6 N_XI803/NET08_XI803/MM6_d N_XI803/QB_XI803/MM6_g N_VDD_XI803/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI803/MM5 N_XI803/Q_XI803/MM5_d N_XI803/QB_XI803/MM5_g N_VDD_XI803/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI803/MM4 N_XI803/QB_XI803/MM4_d N_XI803/Q_XI803/MM4_g N_VDD_XI803/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI802/MM8 N_XI802/NET08_XI802/MM8_d N_RWL<1>_XI802/MM8_g N_RBL<10>_XI802/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI802/MM7 N_XI802/NET08_XI802/MM7_d N_XI802/QB_XI802/MM7_g N_GND_XI802/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI802/MM10 N_WBL<10>_XI802/MM10_d N_WWLB<1>_XI802/MM10_g N_XI802/Q_XI802/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI802/MM11 N_WBLB<10>_XI802/MM11_d N_WWLB<1>_XI802/MM11_g
+ N_XI802/QB_XI802/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI802/MM1 N_XI802/Q_XI802/MM1_d N_XI802/QB_XI802/MM1_g N_GND_XI802/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI802/MM0 N_XI802/QB_XI802/MM0_d N_XI802/Q_XI802/MM0_g N_GND_XI802/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI802/MM9 N_XI802/NET08_XI802/MM9_d N_RWLB<1>_XI802/MM9_g N_RBL<10>_XI802/MM9_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI802/MM6 N_XI802/NET08_XI802/MM6_d N_XI802/QB_XI802/MM6_g N_VDD_XI802/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI802/MM5 N_XI802/Q_XI802/MM5_d N_XI802/QB_XI802/MM5_g N_VDD_XI802/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI802/MM4 N_XI802/QB_XI802/MM4_d N_XI802/Q_XI802/MM4_g N_VDD_XI802/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI807/MM8 N_XI807/NET08_XI807/MM8_d N_RWL<1>_XI807/MM8_g N_RBL<5>_XI807/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI807/MM7 N_XI807/NET08_XI807/MM7_d N_XI807/QB_XI807/MM7_g N_GND_XI807/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI807/MM10 N_WBL<5>_XI807/MM10_d N_WWLB<1>_XI807/MM10_g N_XI807/Q_XI807/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI807/MM11 N_WBLB<5>_XI807/MM11_d N_WWLB<1>_XI807/MM11_g
+ N_XI807/QB_XI807/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI807/MM1 N_XI807/Q_XI807/MM1_d N_XI807/QB_XI807/MM1_g N_GND_XI807/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI807/MM0 N_XI807/QB_XI807/MM0_d N_XI807/Q_XI807/MM0_g N_GND_XI807/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI807/MM9 N_XI807/NET08_XI807/MM9_d N_RWLB<1>_XI807/MM9_g N_RBL<5>_XI807/MM9_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI807/MM6 N_XI807/NET08_XI807/MM6_d N_XI807/QB_XI807/MM6_g N_VDD_XI807/MM6_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI807/MM5 N_XI807/Q_XI807/MM5_d N_XI807/QB_XI807/MM5_g N_VDD_XI807/MM5_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI807/MM4 N_XI807/QB_XI807/MM4_d N_XI807/Q_XI807/MM4_g N_VDD_XI807/MM4_s
+ N_VDD_XI1030/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI835/MM8 N_XI835/NET08_XI835/MM8_d N_RWL<3>_XI835/MM8_g N_RBL<9>_XI835/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI835/MM7 N_XI835/NET08_XI835/MM7_d N_XI835/QB_XI835/MM7_g N_GND_XI835/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI835/MM10 N_WBL<9>_XI835/MM10_d N_WWLB<3>_XI835/MM10_g N_XI835/Q_XI835/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI835/MM11 N_WBLB<9>_XI835/MM11_d N_WWLB<3>_XI835/MM11_g
+ N_XI835/QB_XI835/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI835/MM1 N_XI835/Q_XI835/MM1_d N_XI835/QB_XI835/MM1_g N_GND_XI835/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI835/MM0 N_XI835/QB_XI835/MM0_d N_XI835/Q_XI835/MM0_g N_GND_XI835/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI835/MM9 N_XI835/NET08_XI835/MM9_d N_RWLB<3>_XI835/MM9_g N_RBL<9>_XI835/MM9_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI835/MM6 N_XI835/NET08_XI835/MM6_d N_XI835/QB_XI835/MM6_g N_VDD_XI835/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI835/MM5 N_XI835/Q_XI835/MM5_d N_XI835/QB_XI835/MM5_g N_VDD_XI835/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI835/MM4 N_XI835/QB_XI835/MM4_d N_XI835/Q_XI835/MM4_g N_VDD_XI835/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI834/MM8 N_XI834/NET08_XI834/MM8_d N_RWL<3>_XI834/MM8_g N_RBL<10>_XI834/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI834/MM7 N_XI834/NET08_XI834/MM7_d N_XI834/QB_XI834/MM7_g N_GND_XI834/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI834/MM10 N_WBL<10>_XI834/MM10_d N_WWLB<3>_XI834/MM10_g N_XI834/Q_XI834/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI834/MM11 N_WBLB<10>_XI834/MM11_d N_WWLB<3>_XI834/MM11_g
+ N_XI834/QB_XI834/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI834/MM1 N_XI834/Q_XI834/MM1_d N_XI834/QB_XI834/MM1_g N_GND_XI834/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI834/MM0 N_XI834/QB_XI834/MM0_d N_XI834/Q_XI834/MM0_g N_GND_XI834/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI834/MM9 N_XI834/NET08_XI834/MM9_d N_RWLB<3>_XI834/MM9_g N_RBL<10>_XI834/MM9_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI834/MM6 N_XI834/NET08_XI834/MM6_d N_XI834/QB_XI834/MM6_g N_VDD_XI834/MM6_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI834/MM5 N_XI834/Q_XI834/MM5_d N_XI834/QB_XI834/MM5_g N_VDD_XI834/MM5_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI834/MM4 N_XI834/QB_XI834/MM4_d N_XI834/Q_XI834/MM4_g N_VDD_XI834/MM4_s
+ N_VDD_XI1026/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI833/MM8 N_XI833/NET08_XI833/MM8_d N_RWL<3>_XI833/MM8_g N_RBL<11>_XI833/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI833/MM7 N_XI833/NET08_XI833/MM7_d N_XI833/QB_XI833/MM7_g N_GND_XI833/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI833/MM10 N_WBL<11>_XI833/MM10_d N_WWLB<3>_XI833/MM10_g N_XI833/Q_XI833/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI833/MM11 N_WBLB<11>_XI833/MM11_d N_WWLB<3>_XI833/MM11_g
+ N_XI833/QB_XI833/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI833/MM1 N_XI833/Q_XI833/MM1_d N_XI833/QB_XI833/MM1_g N_GND_XI833/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI833/MM0 N_XI833/QB_XI833/MM0_d N_XI833/Q_XI833/MM0_g N_GND_XI833/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI833/MM9 N_XI833/NET08_XI833/MM9_d N_RWLB<3>_XI833/MM9_g N_RBL<11>_XI833/MM9_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI833/MM6 N_XI833/NET08_XI833/MM6_d N_XI833/QB_XI833/MM6_g N_VDD_XI833/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI833/MM5 N_XI833/Q_XI833/MM5_d N_XI833/QB_XI833/MM5_g N_VDD_XI833/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI833/MM4 N_XI833/QB_XI833/MM4_d N_XI833/Q_XI833/MM4_g N_VDD_XI833/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI832/MM8 N_XI832/NET08_XI832/MM8_d N_RWL<3>_XI832/MM8_g N_RBL<12>_XI832/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI832/MM7 N_XI832/NET08_XI832/MM7_d N_XI832/QB_XI832/MM7_g N_GND_XI832/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI832/MM10 N_WBL<12>_XI832/MM10_d N_WWLB<3>_XI832/MM10_g N_XI832/Q_XI832/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI832/MM11 N_WBLB<12>_XI832/MM11_d N_WWLB<3>_XI832/MM11_g
+ N_XI832/QB_XI832/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI832/MM1 N_XI832/Q_XI832/MM1_d N_XI832/QB_XI832/MM1_g N_GND_XI832/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI832/MM0 N_XI832/QB_XI832/MM0_d N_XI832/Q_XI832/MM0_g N_GND_XI832/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI832/MM9 N_XI832/NET08_XI832/MM9_d N_RWLB<3>_XI832/MM9_g N_RBL<12>_XI832/MM9_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI832/MM6 N_XI832/NET08_XI832/MM6_d N_XI832/QB_XI832/MM6_g N_VDD_XI832/MM6_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI832/MM5 N_XI832/Q_XI832/MM5_d N_XI832/QB_XI832/MM5_g N_VDD_XI832/MM5_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI832/MM4 N_XI832/QB_XI832/MM4_d N_XI832/Q_XI832/MM4_g N_VDD_XI832/MM4_s
+ N_VDD_XI1024/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1022/MM8 N_XI1022/NET08_XI1022/MM8_d N_RWL<15>_XI1022/MM8_g
+ N_RBL<14>_XI1022/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1022/MM7 N_XI1022/NET08_XI1022/MM7_d N_XI1022/QB_XI1022/MM7_g
+ N_GND_XI1022/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1022/MM10 N_WBL<14>_XI1022/MM10_d N_WWLB<15>_XI1022/MM10_g
+ N_XI1022/Q_XI1022/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1022/MM11 N_WBLB<14>_XI1022/MM11_d N_WWLB<15>_XI1022/MM11_g
+ N_XI1022/QB_XI1022/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1022/MM1 N_XI1022/Q_XI1022/MM1_d N_XI1022/QB_XI1022/MM1_g N_GND_XI1022/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1022/MM0 N_XI1022/QB_XI1022/MM0_d N_XI1022/Q_XI1022/MM0_g N_GND_XI1022/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1022/MM9 N_XI1022/NET08_XI1022/MM9_d N_RWLB<15>_XI1022/MM9_g
+ N_RBL<14>_XI1022/MM9_s N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1022/MM6 N_XI1022/NET08_XI1022/MM6_d N_XI1022/QB_XI1022/MM6_g
+ N_VDD_XI1022/MM6_s N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1022/MM5 N_XI1022/Q_XI1022/MM5_d N_XI1022/QB_XI1022/MM5_g N_VDD_XI1022/MM5_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1022/MM4 N_XI1022/QB_XI1022/MM4_d N_XI1022/Q_XI1022/MM4_g N_VDD_XI1022/MM4_s
+ N_VDD_XI1022/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1005/MM8 N_XI1005/NET08_XI1005/MM8_d N_RWL<13>_XI1005/MM8_g
+ N_RBL<15>_XI1005/MM8_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1005/MM7 N_XI1005/NET08_XI1005/MM7_d N_XI1005/QB_XI1005/MM7_g
+ N_GND_XI1005/MM7_s N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1005/MM10 N_WBL<15>_XI1005/MM10_d N_WWLB<13>_XI1005/MM10_g
+ N_XI1005/Q_XI1005/MM10_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1005/MM11 N_WBLB<15>_XI1005/MM11_d N_WWLB<13>_XI1005/MM11_g
+ N_XI1005/QB_XI1005/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI1005/MM1 N_XI1005/Q_XI1005/MM1_d N_XI1005/QB_XI1005/MM1_g N_GND_XI1005/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1005/MM0 N_XI1005/QB_XI1005/MM0_d N_XI1005/Q_XI1005/MM0_g N_GND_XI1005/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI1005/MM9 N_XI1005/NET08_XI1005/MM9_d N_RWLB<13>_XI1005/MM9_g
+ N_RBL<15>_XI1005/MM9_s N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1005/MM6 N_XI1005/NET08_XI1005/MM6_d N_XI1005/QB_XI1005/MM6_g
+ N_VDD_XI1005/MM6_s N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1005/MM5 N_XI1005/Q_XI1005/MM5_d N_XI1005/QB_XI1005/MM5_g N_VDD_XI1005/MM5_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI1005/MM4 N_XI1005/QB_XI1005/MM4_d N_XI1005/Q_XI1005/MM4_g N_VDD_XI1005/MM4_s
+ N_VDD_XI1037/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI789/MM8 N_XI789/NET08_XI789/MM8_d N_RWL<0>_XI789/MM8_g N_RBL<8>_XI789/MM8_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI789/MM7 N_XI789/NET08_XI789/MM7_d N_XI789/QB_XI789/MM7_g N_GND_XI789/MM7_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI789/MM10 N_WBL<8>_XI789/MM10_d N_WWLB<0>_XI789/MM10_g N_XI789/Q_XI789/MM10_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI789/MM11 N_WBLB<8>_XI789/MM11_d N_WWLB<0>_XI789/MM11_g
+ N_XI789/QB_XI789/MM11_s N_GND_XI1037/MM11_b NCH L=6e-08 W=2.4e-07 M=1
mXI789/MM1 N_XI789/Q_XI789/MM1_d N_XI789/QB_XI789/MM1_g N_GND_XI789/MM1_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI789/MM0 N_XI789/QB_XI789/MM0_d N_XI789/Q_XI789/MM0_g N_GND_XI789/MM0_s
+ N_GND_XI1037/MM11_b NCH L=6e-08 W=1.2e-07 M=1
mXI789/MM9 N_XI789/NET08_XI789/MM9_d N_RWLB<0>_XI789/MM9_g N_RBL<8>_XI789/MM9_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI789/MM6 N_XI789/NET08_XI789/MM6_d N_XI789/QB_XI789/MM6_g N_VDD_XI789/MM6_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI789/MM5 N_XI789/Q_XI789/MM5_d N_XI789/QB_XI789/MM5_g N_VDD_XI789/MM5_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
mXI789/MM4 N_XI789/QB_XI789/MM4_d N_XI789/Q_XI789/MM4_g N_VDD_XI789/MM4_s
+ N_VDD_XI1028/MM9_b PCH L=6e-08 W=3.6e-07 M=1
*
.include "/home/wjin/dmtalen/sram/10TSRAM_PEX/16x16_10T_new.pex.netlist.16X16_10T_NEW.pxi"
*
.ends
*
*
